
<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-32.95,39.6893,61.95,-63.2229</PageViewport>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>14.5,-13</position>
<gparam>LABEL_TEXT Go to https://cedar.to/vjyQw7 to download the latest version!</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>14.5,-9.5</position>
<gparam>LABEL_TEXT Error: This file was made with a newer version of Cedar Logic!</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate></page 0>
</circuit>
<throw_away></throw_away>

	<version>2.3.5 | 2018-09-25 23:06:05</version><circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-135.543,38.4453,97.4542,-77.2188</PageViewport>
<gate>
<ID>68</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>-71.5,-173.5</position>
<input>
<ID>ENABLE_0</ID>438 </input>
<input>
<ID>IN_0</ID>259 </input>
<input>
<ID>IN_1</ID>266 </input>
<input>
<ID>IN_10</ID>260 </input>
<input>
<ID>IN_11</ID>261 </input>
<input>
<ID>IN_12</ID>262 </input>
<input>
<ID>IN_13</ID>263 </input>
<input>
<ID>IN_14</ID>264 </input>
<input>
<ID>IN_15</ID>268 </input>
<input>
<ID>IN_2</ID>265 </input>
<input>
<ID>IN_3</ID>255 </input>
<input>
<ID>IN_4</ID>267 </input>
<input>
<ID>IN_5</ID>254 </input>
<input>
<ID>IN_6</ID>253 </input>
<input>
<ID>IN_7</ID>256 </input>
<input>
<ID>IN_8</ID>257 </input>
<input>
<ID>IN_9</ID>258 </input>
<output>
<ID>OUT_0</ID>269 </output>
<output>
<ID>OUT_1</ID>270 </output>
<output>
<ID>OUT_10</ID>284 </output>
<output>
<ID>OUT_11</ID>271 </output>
<output>
<ID>OUT_12</ID>276 </output>
<output>
<ID>OUT_13</ID>272 </output>
<output>
<ID>OUT_14</ID>283 </output>
<output>
<ID>OUT_15</ID>274 </output>
<output>
<ID>OUT_2</ID>278 </output>
<output>
<ID>OUT_3</ID>273 </output>
<output>
<ID>OUT_4</ID>279 </output>
<output>
<ID>OUT_5</ID>277 </output>
<output>
<ID>OUT_6</ID>280 </output>
<output>
<ID>OUT_7</ID>275 </output>
<output>
<ID>OUT_8</ID>281 </output>
<output>
<ID>OUT_9</ID>282 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>4</ID>
<type>AI_RAM_12x16</type>
<position>-26,6</position>
<input>
<ID>ADDRESS_0</ID>6 </input>
<input>
<ID>ADDRESS_1</ID>12 </input>
<input>
<ID>ADDRESS_10</ID>4 </input>
<input>
<ID>ADDRESS_11</ID>2 </input>
<input>
<ID>ADDRESS_2</ID>7 </input>
<input>
<ID>ADDRESS_3</ID>10 </input>
<input>
<ID>ADDRESS_4</ID>5 </input>
<input>
<ID>ADDRESS_5</ID>8 </input>
<input>
<ID>ADDRESS_6</ID>9 </input>
<input>
<ID>ADDRESS_7</ID>11 </input>
<input>
<ID>ADDRESS_8</ID>1 </input>
<input>
<ID>ADDRESS_9</ID>3 </input>
<input>
<ID>DATA_IN_0</ID>18 </input>
<input>
<ID>DATA_IN_1</ID>17 </input>
<input>
<ID>DATA_IN_10</ID>29 </input>
<input>
<ID>DATA_IN_11</ID>23 </input>
<input>
<ID>DATA_IN_12</ID>31 </input>
<input>
<ID>DATA_IN_13</ID>26 </input>
<input>
<ID>DATA_IN_14</ID>25 </input>
<input>
<ID>DATA_IN_15</ID>32 </input>
<input>
<ID>DATA_IN_2</ID>19 </input>
<input>
<ID>DATA_IN_3</ID>27 </input>
<input>
<ID>DATA_IN_4</ID>24 </input>
<input>
<ID>DATA_IN_5</ID>21 </input>
<input>
<ID>DATA_IN_6</ID>22 </input>
<input>
<ID>DATA_IN_7</ID>20 </input>
<input>
<ID>DATA_IN_8</ID>30 </input>
<input>
<ID>DATA_IN_9</ID>28 </input>
<output>
<ID>DATA_OUT_0</ID>18 </output>
<output>
<ID>DATA_OUT_1</ID>17 </output>
<output>
<ID>DATA_OUT_10</ID>29 </output>
<output>
<ID>DATA_OUT_11</ID>23 </output>
<output>
<ID>DATA_OUT_12</ID>31 </output>
<output>
<ID>DATA_OUT_13</ID>26 </output>
<output>
<ID>DATA_OUT_14</ID>25 </output>
<output>
<ID>DATA_OUT_15</ID>32 </output>
<output>
<ID>DATA_OUT_2</ID>19 </output>
<output>
<ID>DATA_OUT_3</ID>27 </output>
<output>
<ID>DATA_OUT_4</ID>24 </output>
<output>
<ID>DATA_OUT_5</ID>21 </output>
<output>
<ID>DATA_OUT_6</ID>22 </output>
<output>
<ID>DATA_OUT_7</ID>20 </output>
<output>
<ID>DATA_OUT_8</ID>30 </output>
<output>
<ID>DATA_OUT_9</ID>28 </output>
<input>
<ID>ENABLE_0</ID>611 </input>
<input>
<ID>write_clock</ID>14 </input>
<input>
<ID>write_enable</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 12</lparam>
<lparam>DATA_BITS 16</lparam>
<lparam>Address:0 16640</lparam>
<lparam>Address:256 8459</lparam>
<lparam>Address:257 12556</lparam>
<lparam>Address:258 8461</lparam>
<lparam>Address:259 12558</lparam>
<lparam>Address:260 30720</lparam>
<lparam>Address:261 37132</lparam>
<lparam>Address:262 24844</lparam>
<lparam>Address:263 24846</lparam>
<lparam>Address:264 16645</lparam>
<lparam>Address:265 12559</lparam>
<lparam>Address:266 28673</lparam>
<lparam>Address:267 336</lparam>
<lparam>Address:268 346</lparam>
<lparam>Address:269 65526</lparam>
<lparam>Address:271 575</lparam>
<lparam>Address:336 25</lparam>
<lparam>Address:337 50</lparam>
<lparam>Address:338 75</lparam>
<lparam>Address:339 100</lparam>
<lparam>Address:340 25</lparam>
<lparam>Address:341 50</lparam>
<lparam>Address:342 75</lparam>
<lparam>Address:343 100</lparam>
<lparam>Address:344 25</lparam>
<lparam>Address:345 50</lparam></gate>
<gate>
<ID>12</ID>
<type>DA_FROM</type>
<position>-14,10.5</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>70</ID>
<type>BX_16X1_BUS_END</type>
<position>-59.5,-173.5</position>
<input>
<ID>Bus_in_0</ID>269 </input>
<input>
<ID>IN_1</ID>270 </input>
<input>
<ID>IN_10</ID>284 </input>
<input>
<ID>IN_11</ID>271 </input>
<input>
<ID>IN_12</ID>276 </input>
<input>
<ID>IN_13</ID>272 </input>
<input>
<ID>IN_14</ID>283 </input>
<input>
<ID>IN_15</ID>274 </input>
<input>
<ID>IN_2</ID>278 </input>
<input>
<ID>IN_3</ID>273 </input>
<input>
<ID>IN_4</ID>279 </input>
<input>
<ID>IN_5</ID>277 </input>
<input>
<ID>IN_6</ID>280 </input>
<input>
<ID>IN_7</ID>275 </input>
<input>
<ID>IN_8</ID>281 </input>
<input>
<ID>IN_9</ID>282 </input>
<input>
<ID>OUT</ID>364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>6</ID>
<type>BX_16X1_BUS_END</type>
<position>-41,8</position>
<input>
<ID>Bus_in_0</ID>6 </input>
<input>
<ID>IN_1</ID>12 </input>
<input>
<ID>IN_10</ID>4 </input>
<input>
<ID>IN_11</ID>2 </input>
<input>
<ID>IN_2</ID>7 </input>
<input>
<ID>IN_3</ID>10 </input>
<input>
<ID>IN_4</ID>5 </input>
<input>
<ID>IN_5</ID>8 </input>
<input>
<ID>IN_6</ID>9 </input>
<input>
<ID>IN_7</ID>11 </input>
<input>
<ID>IN_8</ID>1 </input>
<input>
<ID>IN_9</ID>3 </input>
<input>
<ID>OUT</ID>610 656 689 694 696 735 829 836 860 864 872 873 1001 1002 1003 1016 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>14</ID>
<type>DA_FROM</type>
<position>-15,6.5</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID mem_write</lparam></gate>
<gate>
<ID>17</ID>
<type>BX_16X1_BUS_END</type>
<position>-26,-9</position>
<input>
<ID>Bus_in_0</ID>18 </input>
<input>
<ID>IN_1</ID>17 </input>
<input>
<ID>IN_10</ID>29 </input>
<input>
<ID>IN_11</ID>23 </input>
<input>
<ID>IN_12</ID>31 </input>
<input>
<ID>IN_13</ID>26 </input>
<input>
<ID>IN_14</ID>25 </input>
<input>
<ID>IN_15</ID>32 </input>
<input>
<ID>IN_2</ID>19 </input>
<input>
<ID>IN_3</ID>27 </input>
<input>
<ID>IN_4</ID>24 </input>
<input>
<ID>IN_5</ID>21 </input>
<input>
<ID>IN_6</ID>22 </input>
<input>
<ID>IN_7</ID>20 </input>
<input>
<ID>IN_8</ID>30 </input>
<input>
<ID>IN_9</ID>28 </input>
<input>
<ID>OUT</ID>364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>19</ID>
<type>AI_REGISTER12</type>
<position>-93.5,-35</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>41 </input>
<input>
<ID>IN_10</ID>39 </input>
<input>
<ID>IN_11</ID>35 </input>
<input>
<ID>IN_2</ID>36 </input>
<input>
<ID>IN_3</ID>42 </input>
<input>
<ID>IN_4</ID>40 </input>
<input>
<ID>IN_5</ID>43 </input>
<input>
<ID>IN_6</ID>44 </input>
<input>
<ID>IN_7</ID>34 </input>
<input>
<ID>IN_8</ID>37 </input>
<input>
<ID>IN_9</ID>33 </input>
<output>
<ID>OUT_0</ID>55 </output>
<output>
<ID>OUT_1</ID>49 </output>
<output>
<ID>OUT_10</ID>45 </output>
<output>
<ID>OUT_11</ID>46 </output>
<output>
<ID>OUT_2</ID>50 </output>
<output>
<ID>OUT_3</ID>48 </output>
<output>
<ID>OUT_4</ID>53 </output>
<output>
<ID>OUT_5</ID>47 </output>
<output>
<ID>OUT_6</ID>51 </output>
<output>
<ID>OUT_7</ID>52 </output>
<output>
<ID>OUT_8</ID>56 </output>
<output>
<ID>OUT_9</ID>54 </output>
<input>
<ID>clear</ID>764 </input>
<input>
<ID>clock</ID>416 </input>
<input>
<ID>count_enable</ID>415 </input>
<input>
<ID>load</ID>414 </input>
<gparam>VALUE_BOX -2.4,-0.8,2.4,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 12</lparam>
<lparam>MAX_COUNT 4095</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_LABEL</type>
<position>-104.5,-22</position>
<gparam>LABEL_TEXT Address Register</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>22</ID>
<type>AI_REGISTER12</type>
<position>-93.5,-60</position>
<input>
<ID>IN_0</ID>66 </input>
<input>
<ID>IN_1</ID>63 </input>
<input>
<ID>IN_10</ID>61 </input>
<input>
<ID>IN_11</ID>62 </input>
<input>
<ID>IN_2</ID>64 </input>
<input>
<ID>IN_3</ID>60 </input>
<input>
<ID>IN_4</ID>65 </input>
<input>
<ID>IN_5</ID>58 </input>
<input>
<ID>IN_6</ID>67 </input>
<input>
<ID>IN_7</ID>68 </input>
<input>
<ID>IN_8</ID>59 </input>
<input>
<ID>IN_9</ID>57 </input>
<output>
<ID>OUT_0</ID>81 </output>
<output>
<ID>OUT_1</ID>92 </output>
<output>
<ID>OUT_10</ID>86 </output>
<output>
<ID>OUT_11</ID>91 </output>
<output>
<ID>OUT_2</ID>90 </output>
<output>
<ID>OUT_3</ID>89 </output>
<output>
<ID>OUT_4</ID>84 </output>
<output>
<ID>OUT_5</ID>85 </output>
<output>
<ID>OUT_6</ID>93 </output>
<output>
<ID>OUT_7</ID>88 </output>
<output>
<ID>OUT_8</ID>94 </output>
<output>
<ID>OUT_9</ID>87 </output>
<input>
<ID>clear</ID>824 </input>
<input>
<ID>clock</ID>419 </input>
<input>
<ID>count_enable</ID>418 </input>
<input>
<ID>load</ID>417 </input>
<gparam>VALUE_BOX -2.4,-0.8,2.4,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 267</lparam>
<lparam>INPUT_BITS 12</lparam>
<lparam>MAX_COUNT 4095</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>-105.5,-47.5</position>
<gparam>LABEL_TEXT Program Counter</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>25</ID>
<type>AM_REGISTER16</type>
<position>-93.5,-86.5</position>
<input>
<ID>IN_0</ID>110 </input>
<input>
<ID>IN_1</ID>113 </input>
<input>
<ID>IN_10</ID>122 </input>
<input>
<ID>IN_11</ID>118 </input>
<input>
<ID>IN_12</ID>119 </input>
<input>
<ID>IN_13</ID>123 </input>
<input>
<ID>IN_14</ID>121 </input>
<input>
<ID>IN_15</ID>124 </input>
<input>
<ID>IN_2</ID>109 </input>
<input>
<ID>IN_3</ID>114 </input>
<input>
<ID>IN_4</ID>115 </input>
<input>
<ID>IN_5</ID>116 </input>
<input>
<ID>IN_6</ID>117 </input>
<input>
<ID>IN_7</ID>111 </input>
<input>
<ID>IN_8</ID>112 </input>
<input>
<ID>IN_9</ID>120 </input>
<output>
<ID>OUT_0</ID>129 </output>
<output>
<ID>OUT_1</ID>128 </output>
<output>
<ID>OUT_10</ID>136 </output>
<output>
<ID>OUT_11</ID>125 </output>
<output>
<ID>OUT_12</ID>140 </output>
<output>
<ID>OUT_13</ID>127 </output>
<output>
<ID>OUT_14</ID>137 </output>
<output>
<ID>OUT_15</ID>139 </output>
<output>
<ID>OUT_2</ID>130 </output>
<output>
<ID>OUT_3</ID>131 </output>
<output>
<ID>OUT_4</ID>126 </output>
<output>
<ID>OUT_5</ID>134 </output>
<output>
<ID>OUT_6</ID>135 </output>
<output>
<ID>OUT_7</ID>132 </output>
<output>
<ID>OUT_8</ID>133 </output>
<output>
<ID>OUT_9</ID>138 </output>
<input>
<ID>clock</ID>422 </input>
<input>
<ID>count_enable</ID>421 </input>
<input>
<ID>load</ID>420 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 65536</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>89</ID>
<type>DA_FROM</type>
<position>-110.5,-122.5</position>
<input>
<ID>IN_0</ID>301 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN1</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>-110.5,-72</position>
<gparam>LABEL_TEXT Data Register</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>90</ID>
<type>DA_FROM</type>
<position>-100.5,-121.5</position>
<input>
<ID>IN_0</ID>302 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN2</lparam></gate>
<gate>
<ID>27</ID>
<type>AM_REGISTER16</type>
<position>-93.5,-116</position>
<input>
<ID>IN_0</ID>300 </input>
<input>
<ID>IN_1</ID>301 </input>
<input>
<ID>IN_10</ID>310 </input>
<input>
<ID>IN_11</ID>311 </input>
<input>
<ID>IN_12</ID>312 </input>
<input>
<ID>IN_13</ID>313 </input>
<input>
<ID>IN_14</ID>314 </input>
<input>
<ID>IN_15</ID>315 </input>
<input>
<ID>IN_2</ID>302 </input>
<input>
<ID>IN_3</ID>303 </input>
<input>
<ID>IN_4</ID>304 </input>
<input>
<ID>IN_5</ID>305 </input>
<input>
<ID>IN_6</ID>306 </input>
<input>
<ID>IN_7</ID>307 </input>
<input>
<ID>IN_8</ID>308 </input>
<input>
<ID>IN_9</ID>309 </input>
<output>
<ID>OUT_0</ID>164 </output>
<output>
<ID>OUT_1</ID>161 </output>
<output>
<ID>OUT_10</ID>165 </output>
<output>
<ID>OUT_11</ID>166 </output>
<output>
<ID>OUT_12</ID>158 </output>
<output>
<ID>OUT_13</ID>172 </output>
<output>
<ID>OUT_14</ID>163 </output>
<output>
<ID>OUT_15</ID>170 </output>
<output>
<ID>OUT_2</ID>167 </output>
<output>
<ID>OUT_3</ID>160 </output>
<output>
<ID>OUT_4</ID>159 </output>
<output>
<ID>OUT_5</ID>169 </output>
<output>
<ID>OUT_6</ID>171 </output>
<output>
<ID>OUT_7</ID>162 </output>
<output>
<ID>OUT_8</ID>168 </output>
<output>
<ID>OUT_9</ID>157 </output>
<input>
<ID>clear</ID>426 </input>
<input>
<ID>clock</ID>425 </input>
<input>
<ID>count_enable</ID>424 </input>
<input>
<ID>load</ID>423 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 575</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>91</ID>
<type>DA_FROM</type>
<position>-110.5,-120.5</position>
<input>
<ID>IN_0</ID>303 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN3</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>-108,-104</position>
<gparam>LABEL_TEXT Accumulator</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>92</ID>
<type>DA_FROM</type>
<position>-100.5,-119.5</position>
<input>
<ID>IN_0</ID>304 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN4</lparam></gate>
<gate>
<ID>29</ID>
<type>AM_REGISTER16</type>
<position>-94,-146.5</position>
<input>
<ID>IN_0</ID>190 </input>
<input>
<ID>IN_1</ID>191 </input>
<input>
<ID>IN_10</ID>197 </input>
<input>
<ID>IN_11</ID>200 </input>
<input>
<ID>IN_12</ID>204 </input>
<input>
<ID>IN_13</ID>199 </input>
<input>
<ID>IN_14</ID>203 </input>
<input>
<ID>IN_15</ID>201 </input>
<input>
<ID>IN_2</ID>189 </input>
<input>
<ID>IN_3</ID>192 </input>
<input>
<ID>IN_4</ID>194 </input>
<input>
<ID>IN_5</ID>196 </input>
<input>
<ID>IN_6</ID>195 </input>
<input>
<ID>IN_7</ID>193 </input>
<input>
<ID>IN_8</ID>198 </input>
<input>
<ID>IN_9</ID>202 </input>
<output>
<ID>OUT_0</ID>219 </output>
<output>
<ID>OUT_1</ID>209 </output>
<output>
<ID>OUT_10</ID>218 </output>
<output>
<ID>OUT_11</ID>220 </output>
<output>
<ID>OUT_12</ID>205 </output>
<output>
<ID>OUT_13</ID>207 </output>
<output>
<ID>OUT_14</ID>206 </output>
<output>
<ID>OUT_15</ID>208 </output>
<output>
<ID>OUT_2</ID>210 </output>
<output>
<ID>OUT_3</ID>211 </output>
<output>
<ID>OUT_4</ID>212 </output>
<output>
<ID>OUT_5</ID>213 </output>
<output>
<ID>OUT_6</ID>214 </output>
<output>
<ID>OUT_7</ID>215 </output>
<output>
<ID>OUT_8</ID>216 </output>
<output>
<ID>OUT_9</ID>217 </output>
<input>
<ID>clock</ID>429 </input>
<input>
<ID>load</ID>427 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 28673</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>93</ID>
<type>DA_FROM</type>
<position>-110.5,-118.5</position>
<input>
<ID>IN_0</ID>305 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN5</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>-109,-136</position>
<gparam>LABEL_TEXT Instruction Register</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>94</ID>
<type>DA_FROM</type>
<position>-100.5,-117.5</position>
<input>
<ID>IN_0</ID>306 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN6</lparam></gate>
<gate>
<ID>31</ID>
<type>AM_REGISTER16</type>
<position>-94.5,-173.5</position>
<input>
<ID>IN_0</ID>239 </input>
<input>
<ID>IN_1</ID>238 </input>
<input>
<ID>IN_10</ID>248 </input>
<input>
<ID>IN_11</ID>243 </input>
<input>
<ID>IN_12</ID>251 </input>
<input>
<ID>IN_13</ID>245 </input>
<input>
<ID>IN_14</ID>242 </input>
<input>
<ID>IN_15</ID>247 </input>
<input>
<ID>IN_2</ID>240 </input>
<input>
<ID>IN_3</ID>241 </input>
<input>
<ID>IN_4</ID>237 </input>
<input>
<ID>IN_5</ID>249 </input>
<input>
<ID>IN_6</ID>246 </input>
<input>
<ID>IN_7</ID>250 </input>
<input>
<ID>IN_8</ID>252 </input>
<input>
<ID>IN_9</ID>244 </input>
<output>
<ID>OUT_0</ID>259 </output>
<output>
<ID>OUT_1</ID>266 </output>
<output>
<ID>OUT_10</ID>260 </output>
<output>
<ID>OUT_11</ID>261 </output>
<output>
<ID>OUT_12</ID>262 </output>
<output>
<ID>OUT_13</ID>263 </output>
<output>
<ID>OUT_14</ID>264 </output>
<output>
<ID>OUT_15</ID>268 </output>
<output>
<ID>OUT_2</ID>265 </output>
<output>
<ID>OUT_3</ID>255 </output>
<output>
<ID>OUT_4</ID>267 </output>
<output>
<ID>OUT_5</ID>254 </output>
<output>
<ID>OUT_6</ID>253 </output>
<output>
<ID>OUT_7</ID>256 </output>
<output>
<ID>OUT_8</ID>257 </output>
<output>
<ID>OUT_9</ID>258 </output>
<input>
<ID>clock</ID>432 </input>
<input>
<ID>load</ID>430 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>95</ID>
<type>DA_FROM</type>
<position>-110.5,-116.5</position>
<input>
<ID>IN_0</ID>307 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN7</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>-109,-162.5</position>
<gparam>LABEL_TEXT Temporary Register</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>96</ID>
<type>DA_FROM</type>
<position>-100.5,-115.5</position>
<input>
<ID>IN_0</ID>308 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN8</lparam></gate>
<gate>
<ID>34</ID>
<type>BX_16X1_BUS_END</type>
<position>-102.5,-33</position>
<input>
<ID>Bus_in_0</ID>38 </input>
<input>
<ID>IN_1</ID>41 </input>
<input>
<ID>IN_10</ID>39 </input>
<input>
<ID>IN_11</ID>35 </input>
<input>
<ID>IN_2</ID>36 </input>
<input>
<ID>IN_3</ID>42 </input>
<input>
<ID>IN_4</ID>40 </input>
<input>
<ID>IN_5</ID>43 </input>
<input>
<ID>IN_6</ID>44 </input>
<input>
<ID>IN_7</ID>34 </input>
<input>
<ID>IN_8</ID>37 </input>
<input>
<ID>IN_9</ID>33 </input>
<input>
<ID>OUT</ID>364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>98</ID>
<type>DA_FROM</type>
<position>-100.5,-113.5</position>
<input>
<ID>IN_0</ID>310 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN10</lparam></gate>
<gate>
<ID>38</ID>
<type>BX_16X1_BUS_END</type>
<position>-82,-33</position>
<input>
<ID>Bus_in_0</ID>55 </input>
<input>
<ID>IN_1</ID>49 </input>
<input>
<ID>IN_10</ID>45 </input>
<input>
<ID>IN_11</ID>46 </input>
<input>
<ID>IN_12</ID>1061 </input>
<input>
<ID>IN_13</ID>1061 </input>
<input>
<ID>IN_14</ID>1061 </input>
<input>
<ID>IN_15</ID>1061 </input>
<input>
<ID>IN_2</ID>50 </input>
<input>
<ID>IN_3</ID>48 </input>
<input>
<ID>IN_4</ID>53 </input>
<input>
<ID>IN_5</ID>47 </input>
<input>
<ID>IN_6</ID>51 </input>
<input>
<ID>IN_7</ID>52 </input>
<input>
<ID>IN_8</ID>56 </input>
<input>
<ID>IN_9</ID>54 </input>
<input>
<ID>OUT</ID>610 656 689 694 696 735 829 836 860 864 872 873 1001 1002 1003 1016 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>102</ID>
<type>DA_FROM</type>
<position>-100.5,-109.5</position>
<input>
<ID>IN_0</ID>314 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN14</lparam></gate>
<gate>
<ID>40</ID>
<type>BX_16X1_BUS_END</type>
<position>-103.5,-58</position>
<input>
<ID>Bus_in_0</ID>66 </input>
<input>
<ID>IN_1</ID>63 </input>
<input>
<ID>IN_10</ID>61 </input>
<input>
<ID>IN_11</ID>62 </input>
<input>
<ID>IN_2</ID>64 </input>
<input>
<ID>IN_3</ID>60 </input>
<input>
<ID>IN_4</ID>65 </input>
<input>
<ID>IN_5</ID>58 </input>
<input>
<ID>IN_6</ID>67 </input>
<input>
<ID>IN_7</ID>68 </input>
<input>
<ID>IN_8</ID>59 </input>
<input>
<ID>IN_9</ID>57 </input>
<input>
<ID>OUT</ID>364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>42</ID>
<type>BX_16X1_BUS_END</type>
<position>-75.5,-58</position>
<input>
<ID>Bus_in_0</ID>82 </input>
<input>
<ID>IN_1</ID>83 </input>
<input>
<ID>IN_10</ID>101 </input>
<input>
<ID>IN_11</ID>103 </input>
<input>
<ID>IN_2</ID>108 </input>
<input>
<ID>IN_3</ID>100 </input>
<input>
<ID>IN_4</ID>105 </input>
<input>
<ID>IN_5</ID>102 </input>
<input>
<ID>IN_6</ID>106 </input>
<input>
<ID>IN_7</ID>98 </input>
<input>
<ID>IN_8</ID>99 </input>
<input>
<ID>IN_9</ID>107 </input>
<input>
<ID>OUT</ID>364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>44</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>-82.5,-58</position>
<input>
<ID>ENABLE_0</ID>434 </input>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>92 </input>
<input>
<ID>IN_10</ID>86 </input>
<input>
<ID>IN_11</ID>91 </input>
<input>
<ID>IN_2</ID>90 </input>
<input>
<ID>IN_3</ID>89 </input>
<input>
<ID>IN_4</ID>84 </input>
<input>
<ID>IN_5</ID>85 </input>
<input>
<ID>IN_6</ID>93 </input>
<input>
<ID>IN_7</ID>88 </input>
<input>
<ID>IN_8</ID>94 </input>
<input>
<ID>IN_9</ID>87 </input>
<output>
<ID>OUT_0</ID>82 </output>
<output>
<ID>OUT_1</ID>83 </output>
<output>
<ID>OUT_10</ID>101 </output>
<output>
<ID>OUT_11</ID>103 </output>
<output>
<ID>OUT_2</ID>108 </output>
<output>
<ID>OUT_3</ID>100 </output>
<output>
<ID>OUT_4</ID>105 </output>
<output>
<ID>OUT_5</ID>102 </output>
<output>
<ID>OUT_6</ID>106 </output>
<output>
<ID>OUT_7</ID>98 </output>
<output>
<ID>OUT_8</ID>99 </output>
<output>
<ID>OUT_9</ID>107 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>46</ID>
<type>BX_16X1_BUS_END</type>
<position>-102.5,-86.5</position>
<input>
<ID>Bus_in_0</ID>110 </input>
<input>
<ID>IN_1</ID>113 </input>
<input>
<ID>IN_10</ID>122 </input>
<input>
<ID>IN_11</ID>118 </input>
<input>
<ID>IN_12</ID>119 </input>
<input>
<ID>IN_13</ID>123 </input>
<input>
<ID>IN_14</ID>121 </input>
<input>
<ID>IN_15</ID>124 </input>
<input>
<ID>IN_2</ID>109 </input>
<input>
<ID>IN_3</ID>114 </input>
<input>
<ID>IN_4</ID>115 </input>
<input>
<ID>IN_5</ID>116 </input>
<input>
<ID>IN_6</ID>117 </input>
<input>
<ID>IN_7</ID>111 </input>
<input>
<ID>IN_8</ID>112 </input>
<input>
<ID>IN_9</ID>120 </input>
<input>
<ID>OUT</ID>364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>48</ID>
<type>BX_16X1_BUS_END</type>
<position>-34.5,-86.5</position>
<input>
<ID>Bus_in_0</ID>143 </input>
<input>
<ID>IN_1</ID>144 </input>
<input>
<ID>IN_10</ID>152 </input>
<input>
<ID>IN_11</ID>156 </input>
<input>
<ID>IN_12</ID>543 </input>
<input>
<ID>IN_13</ID>545 </input>
<input>
<ID>IN_14</ID>548 </input>
<input>
<ID>IN_15</ID>550 </input>
<input>
<ID>IN_2</ID>146 </input>
<input>
<ID>IN_3</ID>145 </input>
<input>
<ID>IN_4</ID>147 </input>
<input>
<ID>IN_5</ID>141 </input>
<input>
<ID>IN_6</ID>142 </input>
<input>
<ID>IN_7</ID>154 </input>
<input>
<ID>IN_8</ID>149 </input>
<input>
<ID>IN_9</ID>155 </input>
<input>
<ID>OUT</ID>364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>50</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>-43,-86.5</position>
<input>
<ID>ENABLE_0</ID>435 </input>
<input>
<ID>IN_0</ID>129 </input>
<input>
<ID>IN_1</ID>128 </input>
<input>
<ID>IN_10</ID>136 </input>
<input>
<ID>IN_11</ID>125 </input>
<input>
<ID>IN_12</ID>140 </input>
<input>
<ID>IN_13</ID>127 </input>
<input>
<ID>IN_14</ID>137 </input>
<input>
<ID>IN_15</ID>139 </input>
<input>
<ID>IN_2</ID>130 </input>
<input>
<ID>IN_3</ID>131 </input>
<input>
<ID>IN_4</ID>126 </input>
<input>
<ID>IN_5</ID>134 </input>
<input>
<ID>IN_6</ID>135 </input>
<input>
<ID>IN_7</ID>132 </input>
<input>
<ID>IN_8</ID>133 </input>
<input>
<ID>IN_9</ID>138 </input>
<output>
<ID>OUT_0</ID>143 </output>
<output>
<ID>OUT_1</ID>144 </output>
<output>
<ID>OUT_10</ID>152 </output>
<output>
<ID>OUT_11</ID>156 </output>
<output>
<ID>OUT_12</ID>543 </output>
<output>
<ID>OUT_13</ID>545 </output>
<output>
<ID>OUT_14</ID>548 </output>
<output>
<ID>OUT_15</ID>550 </output>
<output>
<ID>OUT_2</ID>146 </output>
<output>
<ID>OUT_3</ID>145 </output>
<output>
<ID>OUT_4</ID>147 </output>
<output>
<ID>OUT_5</ID>141 </output>
<output>
<ID>OUT_6</ID>142 </output>
<output>
<ID>OUT_7</ID>154 </output>
<output>
<ID>OUT_8</ID>149 </output>
<output>
<ID>OUT_9</ID>155 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>52</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>-47,-116</position>
<input>
<ID>ENABLE_0</ID>436 </input>
<input>
<ID>IN_0</ID>164 </input>
<input>
<ID>IN_1</ID>161 </input>
<input>
<ID>IN_10</ID>165 </input>
<input>
<ID>IN_11</ID>166 </input>
<input>
<ID>IN_12</ID>158 </input>
<input>
<ID>IN_13</ID>172 </input>
<input>
<ID>IN_14</ID>163 </input>
<input>
<ID>IN_15</ID>170 </input>
<input>
<ID>IN_2</ID>167 </input>
<input>
<ID>IN_3</ID>160 </input>
<input>
<ID>IN_4</ID>159 </input>
<input>
<ID>IN_5</ID>169 </input>
<input>
<ID>IN_6</ID>171 </input>
<input>
<ID>IN_7</ID>162 </input>
<input>
<ID>IN_8</ID>168 </input>
<input>
<ID>IN_9</ID>157 </input>
<output>
<ID>OUT_0</ID>182 </output>
<output>
<ID>OUT_1</ID>177 </output>
<output>
<ID>OUT_10</ID>176 </output>
<output>
<ID>OUT_11</ID>174 </output>
<output>
<ID>OUT_12</ID>178 </output>
<output>
<ID>OUT_13</ID>180 </output>
<output>
<ID>OUT_14</ID>181 </output>
<output>
<ID>OUT_15</ID>183 </output>
<output>
<ID>OUT_2</ID>173 </output>
<output>
<ID>OUT_3</ID>188 </output>
<output>
<ID>OUT_4</ID>186 </output>
<output>
<ID>OUT_5</ID>184 </output>
<output>
<ID>OUT_6</ID>179 </output>
<output>
<ID>OUT_7</ID>185 </output>
<output>
<ID>OUT_8</ID>175 </output>
<output>
<ID>OUT_9</ID>187 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>56</ID>
<type>BX_16X1_BUS_END</type>
<position>-34.5,-116</position>
<input>
<ID>Bus_in_0</ID>182 </input>
<input>
<ID>IN_1</ID>177 </input>
<input>
<ID>IN_10</ID>176 </input>
<input>
<ID>IN_11</ID>174 </input>
<input>
<ID>IN_12</ID>178 </input>
<input>
<ID>IN_13</ID>180 </input>
<input>
<ID>IN_14</ID>181 </input>
<input>
<ID>IN_15</ID>183 </input>
<input>
<ID>IN_2</ID>173 </input>
<input>
<ID>IN_3</ID>188 </input>
<input>
<ID>IN_4</ID>186 </input>
<input>
<ID>IN_5</ID>184 </input>
<input>
<ID>IN_6</ID>179 </input>
<input>
<ID>IN_7</ID>185 </input>
<input>
<ID>IN_8</ID>175 </input>
<input>
<ID>IN_9</ID>187 </input>
<input>
<ID>OUT</ID>364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>58</ID>
<type>BX_16X1_BUS_END</type>
<position>-106.5,-146.5</position>
<input>
<ID>Bus_in_0</ID>190 </input>
<input>
<ID>IN_1</ID>191 </input>
<input>
<ID>IN_10</ID>197 </input>
<input>
<ID>IN_11</ID>200 </input>
<input>
<ID>IN_12</ID>204 </input>
<input>
<ID>IN_13</ID>199 </input>
<input>
<ID>IN_14</ID>203 </input>
<input>
<ID>IN_15</ID>201 </input>
<input>
<ID>IN_2</ID>189 </input>
<input>
<ID>IN_3</ID>192 </input>
<input>
<ID>IN_4</ID>194 </input>
<input>
<ID>IN_5</ID>196 </input>
<input>
<ID>IN_6</ID>195 </input>
<input>
<ID>IN_7</ID>193 </input>
<input>
<ID>IN_8</ID>198 </input>
<input>
<ID>IN_9</ID>202 </input>
<input>
<ID>OUT</ID>364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>60</ID>
<type>BX_16X1_BUS_END</type>
<position>-34.5,-146.5</position>
<input>
<ID>Bus_in_0</ID>228 </input>
<input>
<ID>IN_1</ID>232 </input>
<input>
<ID>IN_10</ID>231 </input>
<input>
<ID>IN_11</ID>224 </input>
<input>
<ID>IN_12</ID>225 </input>
<input>
<ID>IN_13</ID>226 </input>
<input>
<ID>IN_14</ID>236 </input>
<input>
<ID>IN_15</ID>235 </input>
<input>
<ID>IN_2</ID>221 </input>
<input>
<ID>IN_3</ID>222 </input>
<input>
<ID>IN_4</ID>227 </input>
<input>
<ID>IN_5</ID>229 </input>
<input>
<ID>IN_6</ID>233 </input>
<input>
<ID>IN_7</ID>234 </input>
<input>
<ID>IN_8</ID>230 </input>
<input>
<ID>IN_9</ID>223 </input>
<input>
<ID>OUT</ID>364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>62</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>-44,-146.5</position>
<input>
<ID>ENABLE_0</ID>437 </input>
<input>
<ID>IN_0</ID>219 </input>
<input>
<ID>IN_1</ID>209 </input>
<input>
<ID>IN_10</ID>218 </input>
<input>
<ID>IN_11</ID>220 </input>
<input>
<ID>IN_12</ID>205 </input>
<input>
<ID>IN_13</ID>207 </input>
<input>
<ID>IN_14</ID>206 </input>
<input>
<ID>IN_15</ID>208 </input>
<input>
<ID>IN_2</ID>210 </input>
<input>
<ID>IN_3</ID>211 </input>
<input>
<ID>IN_4</ID>212 </input>
<input>
<ID>IN_5</ID>213 </input>
<input>
<ID>IN_6</ID>214 </input>
<input>
<ID>IN_7</ID>215 </input>
<input>
<ID>IN_8</ID>216 </input>
<input>
<ID>IN_9</ID>217 </input>
<output>
<ID>OUT_0</ID>228 </output>
<output>
<ID>OUT_1</ID>232 </output>
<output>
<ID>OUT_10</ID>231 </output>
<output>
<ID>OUT_11</ID>224 </output>
<output>
<ID>OUT_12</ID>225 </output>
<output>
<ID>OUT_13</ID>226 </output>
<output>
<ID>OUT_14</ID>236 </output>
<output>
<ID>OUT_15</ID>235 </output>
<output>
<ID>OUT_2</ID>221 </output>
<output>
<ID>OUT_3</ID>222 </output>
<output>
<ID>OUT_4</ID>227 </output>
<output>
<ID>OUT_5</ID>229 </output>
<output>
<ID>OUT_6</ID>233 </output>
<output>
<ID>OUT_7</ID>234 </output>
<output>
<ID>OUT_8</ID>230 </output>
<output>
<ID>OUT_9</ID>223 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>66</ID>
<type>BX_16X1_BUS_END</type>
<position>-107.5,-173.5</position>
<input>
<ID>Bus_in_0</ID>239 </input>
<input>
<ID>IN_1</ID>238 </input>
<input>
<ID>IN_10</ID>248 </input>
<input>
<ID>IN_11</ID>243 </input>
<input>
<ID>IN_12</ID>251 </input>
<input>
<ID>IN_13</ID>245 </input>
<input>
<ID>IN_14</ID>242 </input>
<input>
<ID>IN_15</ID>247 </input>
<input>
<ID>IN_2</ID>240 </input>
<input>
<ID>IN_3</ID>241 </input>
<input>
<ID>IN_4</ID>237 </input>
<input>
<ID>IN_5</ID>249 </input>
<input>
<ID>IN_6</ID>246 </input>
<input>
<ID>IN_7</ID>250 </input>
<input>
<ID>IN_8</ID>252 </input>
<input>
<ID>IN_9</ID>244 </input>
<input>
<ID>OUT</ID>364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>88</ID>
<type>DA_FROM</type>
<position>-100.5,-123.5</position>
<input>
<ID>IN_0</ID>300 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN0</lparam></gate>
<gate>
<ID>97</ID>
<type>DA_FROM</type>
<position>-110.5,-114.5</position>
<input>
<ID>IN_0</ID>309 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN9</lparam></gate>
<gate>
<ID>99</ID>
<type>DA_FROM</type>
<position>-110.5,-112.5</position>
<input>
<ID>IN_0</ID>311 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN11</lparam></gate>
<gate>
<ID>100</ID>
<type>DA_FROM</type>
<position>-100.5,-111.5</position>
<input>
<ID>IN_0</ID>312 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN12</lparam></gate>
<gate>
<ID>101</ID>
<type>DA_FROM</type>
<position>-110.5,-110.5</position>
<input>
<ID>IN_0</ID>313 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN13</lparam></gate>
<gate>
<ID>103</ID>
<type>DA_FROM</type>
<position>-110.5,-108.5</position>
<input>
<ID>IN_0</ID>315 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN15</lparam></gate>
<gate>
<ID>105</ID>
<type>BX_16X1_BUS_END</type>
<position>-61.5,-33</position>
<input>
<ID>Bus_in_0</ID>316 </input>
<input>
<ID>IN_1</ID>317 </input>
<input>
<ID>IN_10</ID>324 </input>
<input>
<ID>IN_11</ID>321 </input>
<input>
<ID>IN_12</ID>1038 </input>
<input>
<ID>IN_13</ID>1039 </input>
<input>
<ID>IN_14</ID>1040 </input>
<input>
<ID>IN_15</ID>1044 </input>
<input>
<ID>IN_2</ID>318 </input>
<input>
<ID>IN_3</ID>319 </input>
<input>
<ID>IN_4</ID>320 </input>
<input>
<ID>IN_5</ID>325 </input>
<input>
<ID>IN_6</ID>329 </input>
<input>
<ID>IN_7</ID>327 </input>
<input>
<ID>IN_8</ID>330 </input>
<input>
<ID>IN_9</ID>326 </input>
<input>
<ID>OUT</ID>610 656 689 694 696 735 829 836 860 864 872 873 1001 1002 1003 1016 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>107</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>-53,-33</position>
<input>
<ID>ENABLE_0</ID>433 </input>
<input>
<ID>IN_0</ID>316 </input>
<input>
<ID>IN_1</ID>317 </input>
<input>
<ID>IN_10</ID>324 </input>
<input>
<ID>IN_11</ID>321 </input>
<input>
<ID>IN_12</ID>1038 </input>
<input>
<ID>IN_13</ID>1039 </input>
<input>
<ID>IN_14</ID>1040 </input>
<input>
<ID>IN_15</ID>1044 </input>
<input>
<ID>IN_2</ID>318 </input>
<input>
<ID>IN_3</ID>319 </input>
<input>
<ID>IN_4</ID>320 </input>
<input>
<ID>IN_5</ID>325 </input>
<input>
<ID>IN_6</ID>329 </input>
<input>
<ID>IN_7</ID>327 </input>
<input>
<ID>IN_8</ID>330 </input>
<input>
<ID>IN_9</ID>326 </input>
<output>
<ID>OUT_0</ID>337 </output>
<output>
<ID>OUT_1</ID>346 </output>
<output>
<ID>OUT_10</ID>340 </output>
<output>
<ID>OUT_11</ID>342 </output>
<output>
<ID>OUT_12</ID>1027 </output>
<output>
<ID>OUT_13</ID>1033 </output>
<output>
<ID>OUT_14</ID>1036 </output>
<output>
<ID>OUT_15</ID>1037 </output>
<output>
<ID>OUT_2</ID>334 </output>
<output>
<ID>OUT_3</ID>335 </output>
<output>
<ID>OUT_4</ID>338 </output>
<output>
<ID>OUT_5</ID>332 </output>
<output>
<ID>OUT_6</ID>336 </output>
<output>
<ID>OUT_7</ID>339 </output>
<output>
<ID>OUT_8</ID>347 </output>
<output>
<ID>OUT_9</ID>341 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>109</ID>
<type>BX_16X1_BUS_END</type>
<position>-40,-33</position>
<input>
<ID>Bus_in_0</ID>337 </input>
<input>
<ID>IN_1</ID>346 </input>
<input>
<ID>IN_10</ID>340 </input>
<input>
<ID>IN_11</ID>342 </input>
<input>
<ID>IN_12</ID>1027 </input>
<input>
<ID>IN_13</ID>1033 </input>
<input>
<ID>IN_14</ID>1036 </input>
<input>
<ID>IN_15</ID>1037 </input>
<input>
<ID>IN_2</ID>334 </input>
<input>
<ID>IN_3</ID>335 </input>
<input>
<ID>IN_4</ID>338 </input>
<input>
<ID>IN_5</ID>332 </input>
<input>
<ID>IN_6</ID>336 </input>
<input>
<ID>IN_7</ID>339 </input>
<input>
<ID>IN_8</ID>347 </input>
<input>
<ID>IN_9</ID>341 </input>
<input>
<ID>OUT</ID>364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>111</ID>
<type>BX_16X1_BUS_END</type>
<position>14.5,-14.5</position>
<input>
<ID>Bus_in_0</ID>410 </input>
<input>
<ID>IN_1</ID>399 </input>
<input>
<ID>IN_10</ID>408 </input>
<input>
<ID>IN_11</ID>396 </input>
<input>
<ID>IN_12</ID>407 </input>
<input>
<ID>IN_13</ID>402 </input>
<input>
<ID>IN_14</ID>403 </input>
<input>
<ID>IN_15</ID>411 </input>
<input>
<ID>IN_2</ID>400 </input>
<input>
<ID>IN_3</ID>409 </input>
<input>
<ID>IN_4</ID>398 </input>
<input>
<ID>IN_5</ID>401 </input>
<input>
<ID>IN_6</ID>397 </input>
<input>
<ID>IN_7</ID>406 </input>
<input>
<ID>IN_8</ID>404 </input>
<input>
<ID>IN_9</ID>405 </input>
<input>
<ID>OUT</ID>364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>113</ID>
<type>AM_REGISTER16</type>
<position>26,-14.5</position>
<input>
<ID>IN_0</ID>410 </input>
<input>
<ID>IN_1</ID>399 </input>
<input>
<ID>IN_10</ID>408 </input>
<input>
<ID>IN_11</ID>396 </input>
<input>
<ID>IN_12</ID>407 </input>
<input>
<ID>IN_13</ID>402 </input>
<input>
<ID>IN_14</ID>403 </input>
<input>
<ID>IN_15</ID>411 </input>
<input>
<ID>IN_2</ID>400 </input>
<input>
<ID>IN_3</ID>409 </input>
<input>
<ID>IN_4</ID>398 </input>
<input>
<ID>IN_5</ID>401 </input>
<input>
<ID>IN_6</ID>397 </input>
<input>
<ID>IN_7</ID>406 </input>
<input>
<ID>IN_8</ID>404 </input>
<input>
<ID>IN_9</ID>405 </input>
<input>
<ID>clock</ID>412 </input>
<input>
<ID>load</ID>413 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>115</ID>
<type>DA_FROM</type>
<position>25,-27</position>
<input>
<ID>IN_0</ID>412 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>117</ID>
<type>DA_FROM</type>
<position>25,-3</position>
<input>
<ID>IN_0</ID>413 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ldOUTR</lparam></gate>
<gate>
<ID>119</ID>
<type>DA_FROM</type>
<position>-96.5,-25</position>
<input>
<ID>IN_0</ID>414 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ldAR</lparam></gate>
<gate>
<ID>121</ID>
<type>DA_FROM</type>
<position>-93.5,-24.5</position>
<input>
<ID>IN_0</ID>415 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID incAR</lparam></gate>
<gate>
<ID>123</ID>
<type>DA_FROM</type>
<position>-94.5,-44.5</position>
<input>
<ID>IN_0</ID>416 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>125</ID>
<type>DA_FROM</type>
<position>-97,-50.5</position>
<input>
<ID>IN_0</ID>417 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ldPC</lparam></gate>
<gate>
<ID>127</ID>
<type>DA_FROM</type>
<position>-91.5,-49.5</position>
<input>
<ID>IN_0</ID>418 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID incPC</lparam></gate>
<gate>
<ID>129</ID>
<type>DA_FROM</type>
<position>-94.5,-69.5</position>
<input>
<ID>IN_0</ID>419 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>131</ID>
<type>DA_FROM</type>
<position>-98,-74.5</position>
<input>
<ID>IN_0</ID>420 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ldDR</lparam></gate>
<gate>
<ID>133</ID>
<type>DA_FROM</type>
<position>-91.5,-74.5</position>
<input>
<ID>IN_0</ID>421 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID incDR</lparam></gate>
<gate>
<ID>135</ID>
<type>DA_FROM</type>
<position>-94.5,-98</position>
<input>
<ID>IN_0</ID>422 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>137</ID>
<type>DA_FROM</type>
<position>-98,-102.5</position>
<input>
<ID>IN_0</ID>423 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ldAC</lparam></gate>
<gate>
<ID>139</ID>
<type>DA_FROM</type>
<position>-89.5,-102.5</position>
<input>
<ID>IN_0</ID>424 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID incAC</lparam></gate>
<gate>
<ID>141</ID>
<type>DA_FROM</type>
<position>-94.5,-127.5</position>
<input>
<ID>IN_0</ID>425 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>143</ID>
<type>DA_FROM</type>
<position>-92.5,-127.5</position>
<input>
<ID>IN_0</ID>426 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID clrAC</lparam></gate>
<gate>
<ID>145</ID>
<type>DA_FROM</type>
<position>-98,-135</position>
<input>
<ID>IN_0</ID>427 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ldIR</lparam></gate>
<gate>
<ID>149</ID>
<type>DA_FROM</type>
<position>-95,-158</position>
<input>
<ID>IN_0</ID>429 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>151</ID>
<type>DA_FROM</type>
<position>-97.5,-162</position>
<input>
<ID>IN_0</ID>430 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ldTR</lparam></gate>
<gate>
<ID>155</ID>
<type>DA_FROM</type>
<position>-95.5,-185</position>
<input>
<ID>IN_0</ID>432 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>157</ID>
<type>DA_FROM</type>
<position>-53,-22</position>
<input>
<ID>IN_0</ID>433 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID busAR</lparam></gate>
<gate>
<ID>159</ID>
<type>DA_FROM</type>
<position>-79,-46.5</position>
<input>
<ID>IN_0</ID>434 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID busPC</lparam></gate>
<gate>
<ID>161</ID>
<type>DA_FROM</type>
<position>-43,-75.5</position>
<input>
<ID>IN_0</ID>435 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID busDR</lparam></gate>
<gate>
<ID>163</ID>
<type>DA_FROM</type>
<position>-47,-105</position>
<input>
<ID>IN_0</ID>436 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID busAC</lparam></gate>
<gate>
<ID>165</ID>
<type>DA_FROM</type>
<position>-44,-135.5</position>
<input>
<ID>IN_0</ID>437 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID busIR</lparam></gate>
<gate>
<ID>167</ID>
<type>DA_FROM</type>
<position>-71.5,-162.5</position>
<input>
<ID>IN_0</ID>438 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID busTR</lparam></gate>
<gate>
<ID>169</ID>
<type>DE_TO</type>
<position>-86.5,-95.5</position>
<input>
<ID>IN_0</ID>129 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr0</lparam></gate>
<gate>
<ID>170</ID>
<type>DE_TO</type>
<position>-86,-97.5</position>
<input>
<ID>IN_0</ID>128 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr1</lparam></gate>
<gate>
<ID>171</ID>
<type>DE_TO</type>
<position>-85.5,-99.5</position>
<input>
<ID>IN_0</ID>130 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr2</lparam></gate>
<gate>
<ID>172</ID>
<type>DE_TO</type>
<position>-85,-101.5</position>
<input>
<ID>IN_0</ID>131 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr3</lparam></gate>
<gate>
<ID>173</ID>
<type>DE_TO</type>
<position>-79.5,-95.5</position>
<input>
<ID>IN_0</ID>126 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr4</lparam></gate>
<gate>
<ID>174</ID>
<type>DE_TO</type>
<position>-79,-97.5</position>
<input>
<ID>IN_0</ID>134 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr5</lparam></gate>
<gate>
<ID>175</ID>
<type>DE_TO</type>
<position>-78.5,-99.5</position>
<input>
<ID>IN_0</ID>135 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr6</lparam></gate>
<gate>
<ID>176</ID>
<type>DE_TO</type>
<position>-78,-101.5</position>
<input>
<ID>IN_0</ID>132 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr7</lparam></gate>
<gate>
<ID>177</ID>
<type>DE_TO</type>
<position>-72.5,-95.5</position>
<input>
<ID>IN_0</ID>133 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr8</lparam></gate>
<gate>
<ID>178</ID>
<type>DE_TO</type>
<position>-72,-97.5</position>
<input>
<ID>IN_0</ID>138 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr9</lparam></gate>
<gate>
<ID>179</ID>
<type>DE_TO</type>
<position>-71.5,-99.5</position>
<input>
<ID>IN_0</ID>136 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr10</lparam></gate>
<gate>
<ID>180</ID>
<type>DE_TO</type>
<position>-71,-101.5</position>
<input>
<ID>IN_0</ID>125 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr11</lparam></gate>
<gate>
<ID>181</ID>
<type>DE_TO</type>
<position>-64.5,-95.5</position>
<input>
<ID>IN_0</ID>140 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr12</lparam></gate>
<gate>
<ID>182</ID>
<type>DE_TO</type>
<position>-64,-97.5</position>
<input>
<ID>IN_0</ID>127 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr13</lparam></gate>
<gate>
<ID>183</ID>
<type>DE_TO</type>
<position>-63.5,-99.5</position>
<input>
<ID>IN_0</ID>137 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr14</lparam></gate>
<gate>
<ID>184</ID>
<type>DE_TO</type>
<position>-63,-101.5</position>
<input>
<ID>IN_0</ID>139 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr15</lparam></gate>
<gate>
<ID>186</ID>
<type>DE_TO</type>
<position>-86.5,-125</position>
<input>
<ID>IN_0</ID>164 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac0</lparam></gate>
<gate>
<ID>188</ID>
<type>DE_TO</type>
<position>-86,-127</position>
<input>
<ID>IN_0</ID>161 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac1</lparam></gate>
<gate>
<ID>189</ID>
<type>DE_TO</type>
<position>-85.5,-129</position>
<input>
<ID>IN_0</ID>167 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac2</lparam></gate>
<gate>
<ID>190</ID>
<type>DE_TO</type>
<position>-85,-131</position>
<input>
<ID>IN_0</ID>160 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac3</lparam></gate>
<gate>
<ID>191</ID>
<type>DE_TO</type>
<position>-79.5,-125</position>
<input>
<ID>IN_0</ID>159 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac4</lparam></gate>
<gate>
<ID>192</ID>
<type>DE_TO</type>
<position>-79,-127</position>
<input>
<ID>IN_0</ID>169 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac5</lparam></gate>
<gate>
<ID>193</ID>
<type>DE_TO</type>
<position>-78.5,-129</position>
<input>
<ID>IN_0</ID>171 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac6</lparam></gate>
<gate>
<ID>194</ID>
<type>DE_TO</type>
<position>-78,-131</position>
<input>
<ID>IN_0</ID>162 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac7</lparam></gate>
<gate>
<ID>195</ID>
<type>DE_TO</type>
<position>-72.5,-125</position>
<input>
<ID>IN_0</ID>168 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac8</lparam></gate>
<gate>
<ID>196</ID>
<type>DE_TO</type>
<position>-72,-127</position>
<input>
<ID>IN_0</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac9</lparam></gate>
<gate>
<ID>197</ID>
<type>DE_TO</type>
<position>-71.5,-129</position>
<input>
<ID>IN_0</ID>165 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac10</lparam></gate>
<gate>
<ID>198</ID>
<type>DE_TO</type>
<position>-71,-131</position>
<input>
<ID>IN_0</ID>166 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac11</lparam></gate>
<gate>
<ID>199</ID>
<type>DE_TO</type>
<position>-64.5,-125</position>
<input>
<ID>IN_0</ID>158 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac12</lparam></gate>
<gate>
<ID>200</ID>
<type>DE_TO</type>
<position>-64,-127</position>
<input>
<ID>IN_0</ID>172 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac13</lparam></gate>
<gate>
<ID>201</ID>
<type>DE_TO</type>
<position>-63.5,-129</position>
<input>
<ID>IN_0</ID>163 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac14</lparam></gate>
<gate>
<ID>202</ID>
<type>DE_TO</type>
<position>-63,-131</position>
<input>
<ID>IN_0</ID>170 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac15</lparam></gate>
<gate>
<ID>203</ID>
<type>DE_TO</type>
<position>-87,-155.5</position>
<input>
<ID>IN_0</ID>219 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir0</lparam></gate>
<gate>
<ID>204</ID>
<type>DE_TO</type>
<position>-86.5,-157.5</position>
<input>
<ID>IN_0</ID>209 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir1</lparam></gate>
<gate>
<ID>205</ID>
<type>DE_TO</type>
<position>-86,-159.5</position>
<input>
<ID>IN_0</ID>210 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir2</lparam></gate>
<gate>
<ID>206</ID>
<type>DE_TO</type>
<position>-85.5,-161.5</position>
<input>
<ID>IN_0</ID>211 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir3</lparam></gate>
<gate>
<ID>207</ID>
<type>DE_TO</type>
<position>-81,-155.5</position>
<input>
<ID>IN_0</ID>212 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir4</lparam></gate>
<gate>
<ID>208</ID>
<type>DE_TO</type>
<position>-80.5,-157.5</position>
<input>
<ID>IN_0</ID>213 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir5</lparam></gate>
<gate>
<ID>209</ID>
<type>DE_TO</type>
<position>-80,-159.5</position>
<input>
<ID>IN_0</ID>214 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir6</lparam></gate>
<gate>
<ID>210</ID>
<type>DE_TO</type>
<position>-79.5,-161.5</position>
<input>
<ID>IN_0</ID>215 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir7</lparam></gate>
<gate>
<ID>211</ID>
<type>DE_TO</type>
<position>-67,-155.5</position>
<input>
<ID>IN_0</ID>216 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir8</lparam></gate>
<gate>
<ID>212</ID>
<type>DE_TO</type>
<position>-66.5,-157.5</position>
<input>
<ID>IN_0</ID>217 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir9</lparam></gate>
<gate>
<ID>213</ID>
<type>DE_TO</type>
<position>-66,-159.5</position>
<input>
<ID>IN_0</ID>218 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir10</lparam></gate>
<gate>
<ID>214</ID>
<type>DE_TO</type>
<position>-65.5,-161.5</position>
<input>
<ID>IN_0</ID>220 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir11</lparam></gate>
<gate>
<ID>215</ID>
<type>DE_TO</type>
<position>-60,-155.5</position>
<input>
<ID>IN_0</ID>205 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir12</lparam></gate>
<gate>
<ID>216</ID>
<type>DE_TO</type>
<position>-59.5,-157.5</position>
<input>
<ID>IN_0</ID>207 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir13</lparam></gate>
<gate>
<ID>217</ID>
<type>DE_TO</type>
<position>-58.5,-159.5</position>
<input>
<ID>IN_0</ID>206 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir14</lparam></gate>
<gate>
<ID>218</ID>
<type>DE_TO</type>
<position>-58,-161.5</position>
<input>
<ID>IN_0</ID>208 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir15</lparam></gate>
<gate>
<ID>291</ID>
<type>DA_FROM</type>
<position>-15,4</position>
<input>
<ID>IN_0</ID>611 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID mem_read</lparam></gate>
<gate>
<ID>556</ID>
<type>DA_FROM</type>
<position>-88.5,-44.5</position>
<input>
<ID>IN_0</ID>764 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID clrAR</lparam></gate>
<gate>
<ID>759</ID>
<type>DA_FROM</type>
<position>-88.5,-70</position>
<input>
<ID>IN_0</ID>824 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID clrPC</lparam></gate>
<gate>
<ID>539</ID>
<type>FF_GND</type>
<position>-87,-24.5</position>
<output>
<ID>OUT_0</ID>1061 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>30 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-26.5,-7,-26.5,-5</points>
<connection>
<GID>4</GID>
<name>DATA_OUT_8</name></connection>
<connection>
<GID>17</GID>
<name>IN_8</name></connection>
<connection>
<GID>4</GID>
<name>DATA_IN_8</name></connection></vsegment></shape></wire>
<wire>
<ID>261 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89.5,-170,-73.5,-170</points>
<connection>
<GID>31</GID>
<name>OUT_11</name></connection>
<connection>
<GID>68</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>14 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-17,7.5,-17,10.5</points>
<connection>
<GID>4</GID>
<name>write_clock</name></connection>
<intersection>10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-17,10.5,-16,10.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>-17 0</intersection></hsegment></shape></wire>
<wire>
<ID>237 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-105.5,-177,-99.5,-177</points>
<connection>
<GID>31</GID>
<name>IN_4</name></connection>
<connection>
<GID>66</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>262 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89.5,-169,-73.5,-169</points>
<connection>
<GID>31</GID>
<name>OUT_12</name></connection>
<connection>
<GID>68</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>29 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28.5,-7,-28.5,-5</points>
<connection>
<GID>4</GID>
<name>DATA_OUT_10</name></connection>
<connection>
<GID>17</GID>
<name>IN_10</name></connection>
<connection>
<GID>4</GID>
<name>DATA_IN_10</name></connection></vsegment></shape></wire>
<wire>
<ID>438 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-71.5,-164.5,-71.5,-164.5</points>
<connection>
<GID>68</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>167</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>259 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89.5,-181,-73.5,-181</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<connection>
<GID>68</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>241 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-105.5,-178,-99.5,-178</points>
<connection>
<GID>31</GID>
<name>IN_3</name></connection>
<connection>
<GID>66</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>266 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89.5,-180,-73.5,-180</points>
<connection>
<GID>31</GID>
<name>OUT_1</name></connection>
<connection>
<GID>68</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>227 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-42,-150,-36.5,-150</points>
<connection>
<GID>60</GID>
<name>IN_4</name></connection>
<connection>
<GID>62</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>260 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89.5,-171,-73.5,-171</points>
<connection>
<GID>31</GID>
<name>OUT_10</name></connection>
<connection>
<GID>68</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>24 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-7,-22.5,-5</points>
<connection>
<GID>4</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>17</GID>
<name>IN_4</name></connection>
<connection>
<GID>4</GID>
<name>DATA_IN_4</name></connection></vsegment></shape></wire>
<wire>
<ID>263 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89.5,-168,-73.5,-168</points>
<connection>
<GID>31</GID>
<name>OUT_13</name></connection>
<connection>
<GID>68</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>247 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-105.5,-166,-99.5,-166</points>
<connection>
<GID>31</GID>
<name>IN_15</name></connection>
<connection>
<GID>66</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>264 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89.5,-167,-73.5,-167</points>
<connection>
<GID>31</GID>
<name>OUT_14</name></connection>
<connection>
<GID>68</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>235 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-42,-139,-36.5,-139</points>
<connection>
<GID>60</GID>
<name>IN_15</name></connection>
<connection>
<GID>62</GID>
<name>OUT_15</name></connection></hsegment></shape></wire>
<wire>
<ID>268 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89.5,-166,-73.5,-166</points>
<connection>
<GID>31</GID>
<name>OUT_15</name></connection>
<connection>
<GID>68</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>265 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89.5,-179,-73.5,-179</points>
<connection>
<GID>31</GID>
<name>OUT_2</name></connection>
<connection>
<GID>68</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>255 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89.5,-178,-73.5,-178</points>
<connection>
<GID>31</GID>
<name>OUT_3</name></connection>
<connection>
<GID>68</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>272 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-69.5,-168,-61.5,-168</points>
<connection>
<GID>68</GID>
<name>OUT_13</name></connection>
<connection>
<GID>70</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>267 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89.5,-177,-73.5,-177</points>
<connection>
<GID>31</GID>
<name>OUT_4</name></connection>
<connection>
<GID>68</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>254 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89.5,-176,-73.5,-176</points>
<connection>
<GID>31</GID>
<name>OUT_5</name></connection>
<connection>
<GID>68</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>253 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89.5,-175,-73.5,-175</points>
<connection>
<GID>31</GID>
<name>OUT_6</name></connection>
<connection>
<GID>68</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>278 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-69.5,-179,-61.5,-179</points>
<connection>
<GID>68</GID>
<name>OUT_2</name></connection>
<connection>
<GID>70</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>239 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-105.5,-181,-99.5,-181</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<connection>
<GID>66</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>256 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89.5,-174,-73.5,-174</points>
<connection>
<GID>31</GID>
<name>OUT_7</name></connection>
<connection>
<GID>68</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>26 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-31.5,-7,-31.5,-5</points>
<connection>
<GID>4</GID>
<name>DATA_OUT_13</name></connection>
<connection>
<GID>17</GID>
<name>IN_13</name></connection>
<connection>
<GID>4</GID>
<name>DATA_IN_13</name></connection></vsegment></shape></wire>
<wire>
<ID>257 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89.5,-173,-73.5,-173</points>
<connection>
<GID>31</GID>
<name>OUT_8</name></connection>
<connection>
<GID>68</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>233 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-42,-148,-36.5,-148</points>
<connection>
<GID>60</GID>
<name>IN_6</name></connection>
<connection>
<GID>62</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>258 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89.5,-172,-73.5,-172</points>
<connection>
<GID>31</GID>
<name>OUT_9</name></connection>
<connection>
<GID>68</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>269 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-69.5,-181,-61.5,-181</points>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection>
<connection>
<GID>70</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>611 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-17,4,-17,5.5</points>
<connection>
<GID>4</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>291</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>245 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-105.5,-168,-99.5,-168</points>
<connection>
<GID>31</GID>
<name>IN_13</name></connection>
<connection>
<GID>66</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>270 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-69.5,-180,-61.5,-180</points>
<connection>
<GID>68</GID>
<name>OUT_1</name></connection>
<connection>
<GID>70</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>251 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-105.5,-169,-99.5,-169</points>
<connection>
<GID>31</GID>
<name>IN_12</name></connection>
<connection>
<GID>66</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>284 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-69.5,-171,-61.5,-171</points>
<connection>
<GID>68</GID>
<name>OUT_10</name></connection>
<connection>
<GID>70</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>399 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-21,21,-21</points>
<connection>
<GID>113</GID>
<name>IN_1</name></connection>
<connection>
<GID>111</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>32 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33.5,-7,-33.5,-5</points>
<connection>
<GID>4</GID>
<name>DATA_OUT_15</name></connection>
<connection>
<GID>17</GID>
<name>IN_15</name></connection>
<connection>
<GID>4</GID>
<name>DATA_IN_15</name></connection></vsegment></shape></wire>
<wire>
<ID>271 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-69.5,-170,-61.5,-170</points>
<connection>
<GID>68</GID>
<name>OUT_11</name></connection>
<connection>
<GID>70</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>243 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-105.5,-170,-99.5,-170</points>
<connection>
<GID>31</GID>
<name>IN_11</name></connection>
<connection>
<GID>66</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>276 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-69.5,-169,-61.5,-169</points>
<connection>
<GID>68</GID>
<name>OUT_12</name></connection>
<connection>
<GID>70</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>283 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-69.5,-167,-61.5,-167</points>
<connection>
<GID>68</GID>
<name>OUT_14</name></connection>
<connection>
<GID>70</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>249 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-105.5,-176,-99.5,-176</points>
<connection>
<GID>31</GID>
<name>IN_5</name></connection>
<connection>
<GID>66</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>274 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-69.5,-166,-61.5,-166</points>
<connection>
<GID>68</GID>
<name>OUT_15</name></connection>
<connection>
<GID>70</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>273 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-69.5,-178,-61.5,-178</points>
<connection>
<GID>68</GID>
<name>OUT_3</name></connection>
<connection>
<GID>70</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>279 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-69.5,-177,-61.5,-177</points>
<connection>
<GID>68</GID>
<name>OUT_4</name></connection>
<connection>
<GID>70</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>277 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-69.5,-176,-61.5,-176</points>
<connection>
<GID>68</GID>
<name>OUT_5</name></connection>
<connection>
<GID>70</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>7 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-39,2.5,-35,2.5</points>
<connection>
<GID>6</GID>
<name>IN_2</name></connection>
<connection>
<GID>4</GID>
<name>ADDRESS_2</name></connection></hsegment></shape></wire>
<wire>
<ID>135 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-88,-45,-88</points>
<connection>
<GID>25</GID>
<name>OUT_6</name></connection>
<connection>
<GID>50</GID>
<name>IN_6</name></connection>
<intersection>-80.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-80.5,-99.5,-80.5,-88</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>-88 1</intersection></vsegment></shape></wire>
<wire>
<ID>280 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-69.5,-175,-61.5,-175</points>
<connection>
<GID>68</GID>
<name>OUT_6</name></connection>
<connection>
<GID>70</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>275 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-69.5,-174,-61.5,-174</points>
<connection>
<GID>68</GID>
<name>OUT_7</name></connection>
<connection>
<GID>70</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>281 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-69.5,-173,-61.5,-173</points>
<connection>
<GID>68</GID>
<name>OUT_8</name></connection>
<connection>
<GID>70</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>1 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-39,8.5,-35,8.5</points>
<connection>
<GID>6</GID>
<name>IN_8</name></connection>
<connection>
<GID>4</GID>
<name>ADDRESS_8</name></connection></hsegment></shape></wire>
<wire>
<ID>129 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-94,-45,-94</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>-88.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-88.5,-95.5,-88.5,-94</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<intersection>-94 1</intersection></vsegment></shape></wire>
<wire>
<ID>282 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-69.5,-172,-61.5,-172</points>
<connection>
<GID>68</GID>
<name>OUT_9</name></connection>
<connection>
<GID>70</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>6 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-39,0.5,-35,0.5</points>
<connection>
<GID>6</GID>
<name>Bus_in_0</name></connection>
<connection>
<GID>4</GID>
<name>ADDRESS_0</name></connection></hsegment></shape></wire>
<wire>
<ID>12 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-39,1.5,-35,1.5</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<connection>
<GID>4</GID>
<name>ADDRESS_1</name></connection></hsegment></shape></wire>
<wire>
<ID>4 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-39,10.5,-35,10.5</points>
<connection>
<GID>6</GID>
<name>IN_10</name></connection>
<connection>
<GID>4</GID>
<name>ADDRESS_10</name></connection></hsegment></shape></wire>
<wire>
<ID>2 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-39,11.5,-35,11.5</points>
<connection>
<GID>6</GID>
<name>IN_11</name></connection>
<connection>
<GID>4</GID>
<name>ADDRESS_11</name></connection></hsegment></shape></wire>
<wire>
<ID>10 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-39,3.5,-35,3.5</points>
<connection>
<GID>6</GID>
<name>IN_3</name></connection>
<connection>
<GID>4</GID>
<name>ADDRESS_3</name></connection></hsegment></shape></wire>
<wire>
<ID>5 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-39,4.5,-35,4.5</points>
<connection>
<GID>6</GID>
<name>IN_4</name></connection>
<connection>
<GID>4</GID>
<name>ADDRESS_4</name></connection></hsegment></shape></wire>
<wire>
<ID>8 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-39,5.5,-35,5.5</points>
<connection>
<GID>6</GID>
<name>IN_5</name></connection>
<connection>
<GID>4</GID>
<name>ADDRESS_5</name></connection></hsegment></shape></wire>
<wire>
<ID>9 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-39,6.5,-35,6.5</points>
<connection>
<GID>6</GID>
<name>IN_6</name></connection>
<connection>
<GID>4</GID>
<name>ADDRESS_6</name></connection></hsegment></shape></wire>
<wire>
<ID>203 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-104.5,-140,-99,-140</points>
<connection>
<GID>29</GID>
<name>IN_14</name></connection>
<connection>
<GID>58</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-122.5,-189,-122.5,-14.5</points>
<intersection>-189 4</intersection>
<intersection>-173.5 22</intersection>
<intersection>-146.5 8</intersection>
<intersection>-86.5 6</intersection>
<intersection>-58 37</intersection>
<intersection>-33 1</intersection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-122.5,-33,-104.5,-33</points>
<connection>
<GID>34</GID>
<name>OUT</name></connection>
<intersection>-122.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-122.5,-14.5,12.5,-14.5</points>
<connection>
<GID>111</GID>
<name>OUT</name></connection>
<intersection>-122.5 0</intersection>
<intersection>-26 14</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-122.5,-189,-26,-189</points>
<intersection>-122.5 0</intersection>
<intersection>-26 14</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-122.5,-86.5,-104.5,-86.5</points>
<connection>
<GID>46</GID>
<name>OUT</name></connection>
<intersection>-122.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-122.5,-146.5,-108.5,-146.5</points>
<connection>
<GID>58</GID>
<name>OUT</name></connection>
<intersection>-122.5 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-26,-189,-26,-11</points>
<connection>
<GID>17</GID>
<name>OUT</name></connection>
<intersection>-189 4</intersection>
<intersection>-173.5 21</intersection>
<intersection>-146.5 24</intersection>
<intersection>-116 26</intersection>
<intersection>-86.5 28</intersection>
<intersection>-58 36</intersection>
<intersection>-33 32</intersection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>-57.5,-173.5,-26,-173.5</points>
<connection>
<GID>70</GID>
<name>OUT</name></connection>
<intersection>-26 14</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>-122.5,-173.5,-109.5,-173.5</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<intersection>-122.5 0</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>-32.5,-146.5,-26,-146.5</points>
<connection>
<GID>60</GID>
<name>OUT</name></connection>
<intersection>-26 14</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>-32.5,-116,-26,-116</points>
<connection>
<GID>56</GID>
<name>OUT</name></connection>
<intersection>-26 14</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>-32.5,-86.5,-26,-86.5</points>
<connection>
<GID>48</GID>
<name>OUT</name></connection>
<intersection>-26 14</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>-38,-33,-26,-33</points>
<connection>
<GID>109</GID>
<name>OUT</name></connection>
<intersection>-26 14</intersection></hsegment>
<hsegment>
<ID>36</ID>
<points>-73.5,-58,-26,-58</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<intersection>-26 14</intersection></hsegment>
<hsegment>
<ID>37</ID>
<points>-122.5,-58,-105.5,-58</points>
<connection>
<GID>40</GID>
<name>OUT</name></connection>
<intersection>-122.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-39,7.5,-35,7.5</points>
<connection>
<GID>6</GID>
<name>IN_7</name></connection>
<connection>
<GID>4</GID>
<name>ADDRESS_7</name></connection></hsegment></shape></wire>
<wire>
<ID>3 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-39,9.5,-35,9.5</points>
<connection>
<GID>6</GID>
<name>IN_9</name></connection>
<connection>
<GID>4</GID>
<name>ADDRESS_9</name></connection></hsegment></shape></wire>
<wire>
<ID>18 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-18.5,-7,-18.5,-5</points>
<connection>
<GID>4</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>17</GID>
<name>Bus_in_0</name></connection>
<connection>
<GID>4</GID>
<name>DATA_IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>17 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-19.5,-7,-19.5,-5</points>
<connection>
<GID>4</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<connection>
<GID>4</GID>
<name>DATA_IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>23 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29.5,-7,-29.5,-5</points>
<connection>
<GID>4</GID>
<name>DATA_OUT_11</name></connection>
<connection>
<GID>17</GID>
<name>IN_11</name></connection>
<connection>
<GID>4</GID>
<name>DATA_IN_11</name></connection></vsegment></shape></wire>
<wire>
<ID>31 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30.5,-7,-30.5,-5</points>
<connection>
<GID>4</GID>
<name>DATA_OUT_12</name></connection>
<connection>
<GID>17</GID>
<name>IN_12</name></connection>
<connection>
<GID>4</GID>
<name>DATA_IN_12</name></connection></vsegment></shape></wire>
<wire>
<ID>25 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32.5,-7,-32.5,-5</points>
<connection>
<GID>4</GID>
<name>DATA_OUT_14</name></connection>
<connection>
<GID>17</GID>
<name>IN_14</name></connection>
<connection>
<GID>4</GID>
<name>DATA_IN_14</name></connection></vsegment></shape></wire>
<wire>
<ID>19 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20.5,-7,-20.5,-5</points>
<connection>
<GID>4</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>17</GID>
<name>IN_2</name></connection>
<connection>
<GID>4</GID>
<name>DATA_IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>27 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-21.5,-7,-21.5,-5</points>
<connection>
<GID>4</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>17</GID>
<name>IN_3</name></connection>
<connection>
<GID>4</GID>
<name>DATA_IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>21 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23.5,-7,-23.5,-5</points>
<connection>
<GID>4</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>17</GID>
<name>IN_5</name></connection>
<connection>
<GID>4</GID>
<name>DATA_IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>22 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-24.5,-7,-24.5,-5</points>
<connection>
<GID>4</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>17</GID>
<name>IN_6</name></connection>
<connection>
<GID>4</GID>
<name>DATA_IN_6</name></connection></vsegment></shape></wire>
<wire>
<ID>20 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25.5,-7,-25.5,-5</points>
<connection>
<GID>4</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>17</GID>
<name>IN_7</name></connection>
<connection>
<GID>4</GID>
<name>DATA_IN_7</name></connection></vsegment></shape></wire>
<wire>
<ID>28 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-27.5,-7,-27.5,-5</points>
<connection>
<GID>4</GID>
<name>DATA_OUT_9</name></connection>
<connection>
<GID>17</GID>
<name>IN_9</name></connection>
<connection>
<GID>4</GID>
<name>DATA_IN_9</name></connection></vsegment></shape></wire>
<wire>
<ID>15 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-17,6.5,-17,6.5</points>
<connection>
<GID>4</GID>
<name>write_enable</name></connection>
<connection>
<GID>14</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>213 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89,-149,-46,-149</points>
<connection>
<GID>29</GID>
<name>OUT_5</name></connection>
<connection>
<GID>62</GID>
<name>IN_5</name></connection>
<intersection>-82.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-82.5,-157.5,-82.5,-149</points>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<intersection>-149 1</intersection></vsegment></shape></wire>
<wire>
<ID>223 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-42,-145,-36.5,-145</points>
<connection>
<GID>60</GID>
<name>IN_9</name></connection>
<connection>
<GID>62</GID>
<name>OUT_9</name></connection></hsegment></shape></wire>
<wire>
<ID>545 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41,-81,-36.5,-81</points>
<connection>
<GID>48</GID>
<name>IN_13</name></connection>
<connection>
<GID>50</GID>
<name>OUT_13</name></connection></hsegment></shape></wire>
<wire>
<ID>217 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89,-145,-46,-145</points>
<connection>
<GID>29</GID>
<name>OUT_9</name></connection>
<connection>
<GID>62</GID>
<name>IN_9</name></connection>
<intersection>-68.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-68.5,-157.5,-68.5,-145</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>-145 1</intersection></vsegment></shape></wire>
<wire>
<ID>211 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89,-151,-46,-151</points>
<connection>
<GID>29</GID>
<name>OUT_3</name></connection>
<connection>
<GID>62</GID>
<name>IN_3</name></connection>
<intersection>-87.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-87.5,-161.5,-87.5,-151</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<intersection>-151 1</intersection></vsegment></shape></wire>
<wire>
<ID>221 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-42,-152,-36.5,-152</points>
<connection>
<GID>60</GID>
<name>IN_2</name></connection>
<connection>
<GID>62</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>231 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-42,-144,-36.5,-144</points>
<connection>
<GID>60</GID>
<name>IN_10</name></connection>
<connection>
<GID>62</GID>
<name>OUT_10</name></connection></hsegment></shape></wire>
<wire>
<ID>225 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-42,-142,-36.5,-142</points>
<connection>
<GID>60</GID>
<name>IN_12</name></connection>
<connection>
<GID>62</GID>
<name>OUT_12</name></connection></hsegment></shape></wire>
<wire>
<ID>610 656 689 694 696 735 829 836 860 864 872 873 1001 1002 1003 1016 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-80,-33,-63.5,-33</points>
<connection>
<GID>105</GID>
<name>OUT</name></connection>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<intersection>-72.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-72.5,-33,-72.5,8</points>
<intersection>-33 1</intersection>
<intersection>8 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-72.5,8,-43,8</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>-72.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>321 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-59.5,-29.5,-55,-29.5</points>
<connection>
<GID>105</GID>
<name>IN_11</name></connection>
<connection>
<GID>107</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>33 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100.5,-31.5,-98.5,-31.5</points>
<connection>
<GID>19</GID>
<name>IN_9</name></connection>
<connection>
<GID>34</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>117 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100.5,-88,-98.5,-88</points>
<connection>
<GID>25</GID>
<name>IN_6</name></connection>
<connection>
<GID>46</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>184 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-45,-118.5,-36.5,-118.5</points>
<connection>
<GID>52</GID>
<name>OUT_5</name></connection>
<connection>
<GID>56</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>317 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-59.5,-39.5,-55,-39.5</points>
<connection>
<GID>105</GID>
<name>IN_1</name></connection>
<connection>
<GID>107</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>169 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-118.5,-49,-118.5</points>
<connection>
<GID>52</GID>
<name>IN_5</name></connection>
<connection>
<GID>27</GID>
<name>OUT_5</name></connection>
<intersection>-81 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-81,-127,-81,-118.5</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>-118.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>397 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-16,21,-16</points>
<connection>
<GID>113</GID>
<name>IN_6</name></connection>
<connection>
<GID>111</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>38 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100.5,-40.5,-98.5,-40.5</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<connection>
<GID>34</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>41 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100.5,-39.5,-98.5,-39.5</points>
<connection>
<GID>19</GID>
<name>IN_1</name></connection>
<connection>
<GID>34</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>39 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100.5,-30.5,-98.5,-30.5</points>
<connection>
<GID>19</GID>
<name>IN_10</name></connection>
<connection>
<GID>34</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>35 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100.5,-29.5,-98.5,-29.5</points>
<connection>
<GID>19</GID>
<name>IN_11</name></connection>
<connection>
<GID>34</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>36 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100.5,-38.5,-98.5,-38.5</points>
<connection>
<GID>19</GID>
<name>IN_2</name></connection>
<connection>
<GID>34</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>401 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-17,21,-17</points>
<connection>
<GID>113</GID>
<name>IN_5</name></connection>
<connection>
<GID>111</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>42 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100.5,-37.5,-98.5,-37.5</points>
<connection>
<GID>19</GID>
<name>IN_3</name></connection>
<connection>
<GID>34</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>407 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-10,21,-10</points>
<connection>
<GID>113</GID>
<name>IN_12</name></connection>
<connection>
<GID>111</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>40 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100.5,-36.5,-98.5,-36.5</points>
<connection>
<GID>19</GID>
<name>IN_4</name></connection>
<connection>
<GID>34</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>43 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100.5,-35.5,-98.5,-35.5</points>
<connection>
<GID>19</GID>
<name>IN_5</name></connection>
<connection>
<GID>34</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>44 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100.5,-34.5,-98.5,-34.5</points>
<connection>
<GID>19</GID>
<name>IN_6</name></connection>
<connection>
<GID>34</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>34 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100.5,-33.5,-98.5,-33.5</points>
<connection>
<GID>19</GID>
<name>IN_7</name></connection>
<connection>
<GID>34</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>37 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100.5,-32.5,-98.5,-32.5</points>
<connection>
<GID>19</GID>
<name>IN_8</name></connection>
<connection>
<GID>34</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>429 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-95,-156,-95,-156</points>
<connection>
<GID>29</GID>
<name>clock</name></connection>
<connection>
<GID>149</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>764 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-92.5,-42.5,-88.5,-42.5</points>
<connection>
<GID>556</GID>
<name>IN_0</name></connection>
<connection>
<GID>19</GID>
<name>clear</name></connection></hsegment></shape></wire>
<wire>
<ID>416 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-94.5,-42.5,-94.5,-42.5</points>
<connection>
<GID>19</GID>
<name>clock</name></connection>
<connection>
<GID>123</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>48 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-37.5,-84,-37.5</points>
<connection>
<GID>19</GID>
<name>OUT_3</name></connection>
<connection>
<GID>38</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>415 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-93.5,-27.5,-93.5,-26.5</points>
<connection>
<GID>19</GID>
<name>count_enable</name></connection>
<connection>
<GID>121</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>414 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-96.5,-27.5,-96.5,-27</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-96.5,-27.5,-94.5,-27.5</points>
<connection>
<GID>19</GID>
<name>load</name></connection>
<intersection>-96.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>55 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-40.5,-84,-40.5</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<connection>
<GID>38</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>49 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-39.5,-84,-39.5</points>
<connection>
<GID>19</GID>
<name>OUT_1</name></connection>
<connection>
<GID>38</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>45 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-30.5,-84,-30.5</points>
<connection>
<GID>19</GID>
<name>OUT_10</name></connection>
<connection>
<GID>38</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>405 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-13,21,-13</points>
<connection>
<GID>113</GID>
<name>IN_9</name></connection>
<connection>
<GID>111</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>46 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-29.5,-84,-29.5</points>
<connection>
<GID>19</GID>
<name>OUT_11</name></connection>
<connection>
<GID>38</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>409 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-19,21,-19</points>
<connection>
<GID>113</GID>
<name>IN_3</name></connection>
<connection>
<GID>111</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>50 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-38.5,-84,-38.5</points>
<connection>
<GID>19</GID>
<name>OUT_2</name></connection>
<connection>
<GID>38</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>53 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-36.5,-84,-36.5</points>
<connection>
<GID>19</GID>
<name>OUT_4</name></connection>
<connection>
<GID>38</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>47 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-35.5,-84,-35.5</points>
<connection>
<GID>19</GID>
<name>OUT_5</name></connection>
<connection>
<GID>38</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>51 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-34.5,-84,-34.5</points>
<connection>
<GID>19</GID>
<name>OUT_6</name></connection>
<connection>
<GID>38</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>403 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-8,21,-8</points>
<connection>
<GID>113</GID>
<name>IN_14</name></connection>
<connection>
<GID>111</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>52 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-33.5,-84,-33.5</points>
<connection>
<GID>19</GID>
<name>OUT_7</name></connection>
<connection>
<GID>38</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>423 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-98,-106.5,-98,-104.5</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<intersection>-106.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-98,-106.5,-94.5,-106.5</points>
<connection>
<GID>27</GID>
<name>load</name></connection>
<intersection>-98 0</intersection></hsegment></shape></wire>
<wire>
<ID>56 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-32.5,-84,-32.5</points>
<connection>
<GID>19</GID>
<name>OUT_8</name></connection>
<connection>
<GID>38</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>413 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-5,25,-5</points>
<connection>
<GID>113</GID>
<name>load</name></connection>
<connection>
<GID>117</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>54 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-31.5,-84,-31.5</points>
<connection>
<GID>19</GID>
<name>OUT_9</name></connection>
<connection>
<GID>38</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>66 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-101.5,-65.5,-98.5,-65.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<connection>
<GID>40</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>63 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-101.5,-64.5,-98.5,-64.5</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<connection>
<GID>40</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>61 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-101.5,-55.5,-98.5,-55.5</points>
<connection>
<GID>22</GID>
<name>IN_10</name></connection>
<connection>
<GID>40</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>421 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-93.5,-77,-91.5,-77</points>
<connection>
<GID>25</GID>
<name>count_enable</name></connection>
<intersection>-91.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-91.5,-77,-91.5,-76.5</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<intersection>-77 1</intersection></vsegment></shape></wire>
<wire>
<ID>62 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-101.5,-54.5,-98.5,-54.5</points>
<connection>
<GID>22</GID>
<name>IN_11</name></connection>
<connection>
<GID>40</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>64 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-101.5,-63.5,-98.5,-63.5</points>
<connection>
<GID>22</GID>
<name>IN_2</name></connection>
<connection>
<GID>40</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>411 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-7,21,-7</points>
<connection>
<GID>113</GID>
<name>IN_15</name></connection>
<connection>
<GID>111</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>60 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-101.5,-62.5,-98.5,-62.5</points>
<connection>
<GID>22</GID>
<name>IN_3</name></connection>
<connection>
<GID>40</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>65 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-101.5,-61.5,-98.5,-61.5</points>
<connection>
<GID>22</GID>
<name>IN_4</name></connection>
<connection>
<GID>40</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>417 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-97,-52.5,-94.5,-52.5</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<connection>
<GID>22</GID>
<name>load</name></connection></hsegment></shape></wire>
<wire>
<ID>58 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-101.5,-60.5,-98.5,-60.5</points>
<connection>
<GID>22</GID>
<name>IN_5</name></connection>
<connection>
<GID>40</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>67 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-101.5,-59.5,-98.5,-59.5</points>
<connection>
<GID>22</GID>
<name>IN_6</name></connection>
<connection>
<GID>40</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>68 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-101.5,-58.5,-98.5,-58.5</points>
<connection>
<GID>22</GID>
<name>IN_7</name></connection>
<connection>
<GID>40</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>59 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-101.5,-57.5,-98.5,-57.5</points>
<connection>
<GID>22</GID>
<name>IN_8</name></connection>
<connection>
<GID>40</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>57 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-101.5,-56.5,-98.5,-56.5</points>
<connection>
<GID>22</GID>
<name>IN_9</name></connection>
<connection>
<GID>40</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>824 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-88.5,-68,-88.5,-67.5</points>
<connection>
<GID>759</GID>
<name>IN_0</name></connection>
<intersection>-67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-92.5,-67.5,-88.5,-67.5</points>
<connection>
<GID>22</GID>
<name>clear</name></connection>
<intersection>-88.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>419 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-94.5,-67.5,-94.5,-67.5</points>
<connection>
<GID>22</GID>
<name>clock</name></connection>
<connection>
<GID>129</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>418 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-91.5,-52.5,-91.5,-51.5</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-93.5,-52.5,-91.5,-52.5</points>
<connection>
<GID>22</GID>
<name>count_enable</name></connection>
<intersection>-91.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>81 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-88.5,-65.5,-84.5,-65.5</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<connection>
<GID>44</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>92 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-64.5,-84.5,-64.5</points>
<connection>
<GID>22</GID>
<name>OUT_1</name></connection>
<connection>
<GID>44</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>86 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-55.5,-84.5,-55.5</points>
<connection>
<GID>22</GID>
<name>OUT_10</name></connection>
<connection>
<GID>44</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>91 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-54.5,-84.5,-54.5</points>
<connection>
<GID>22</GID>
<name>OUT_11</name></connection>
<connection>
<GID>44</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>90 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-63.5,-84.5,-63.5</points>
<connection>
<GID>22</GID>
<name>OUT_2</name></connection>
<connection>
<GID>44</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>89 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-62.5,-84.5,-62.5</points>
<connection>
<GID>22</GID>
<name>OUT_3</name></connection>
<connection>
<GID>44</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>84 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-61.5,-84.5,-61.5</points>
<connection>
<GID>22</GID>
<name>OUT_4</name></connection>
<connection>
<GID>44</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>85 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-60.5,-84.5,-60.5</points>
<connection>
<GID>22</GID>
<name>OUT_5</name></connection>
<connection>
<GID>44</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>93 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-59.5,-84.5,-59.5</points>
<connection>
<GID>22</GID>
<name>OUT_6</name></connection>
<connection>
<GID>44</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>88 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-58.5,-84.5,-58.5</points>
<connection>
<GID>22</GID>
<name>OUT_7</name></connection>
<connection>
<GID>44</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>94 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-57.5,-84.5,-57.5</points>
<connection>
<GID>22</GID>
<name>OUT_8</name></connection>
<connection>
<GID>44</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>87 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-56.5,-84.5,-56.5</points>
<connection>
<GID>22</GID>
<name>OUT_9</name></connection>
<connection>
<GID>44</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>301 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-108.5,-122.5,-98.5,-122.5</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<connection>
<GID>27</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>110 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100.5,-94,-98.5,-94</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<connection>
<GID>46</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>113 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100.5,-93,-98.5,-93</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<connection>
<GID>46</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>122 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100.5,-84,-98.5,-84</points>
<connection>
<GID>25</GID>
<name>IN_10</name></connection>
<connection>
<GID>46</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>118 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100.5,-83,-98.5,-83</points>
<connection>
<GID>25</GID>
<name>IN_11</name></connection>
<connection>
<GID>46</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>119 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100.5,-82,-98.5,-82</points>
<connection>
<GID>25</GID>
<name>IN_12</name></connection>
<connection>
<GID>46</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>123 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100.5,-81,-98.5,-81</points>
<connection>
<GID>25</GID>
<name>IN_13</name></connection>
<connection>
<GID>46</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>121 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100.5,-80,-98.5,-80</points>
<connection>
<GID>25</GID>
<name>IN_14</name></connection>
<connection>
<GID>46</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>124 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100.5,-79,-98.5,-79</points>
<connection>
<GID>25</GID>
<name>IN_15</name></connection>
<connection>
<GID>46</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>109 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100.5,-92,-98.5,-92</points>
<connection>
<GID>25</GID>
<name>IN_2</name></connection>
<connection>
<GID>46</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>114 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100.5,-91,-98.5,-91</points>
<connection>
<GID>25</GID>
<name>IN_3</name></connection>
<connection>
<GID>46</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>115 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100.5,-90,-98.5,-90</points>
<connection>
<GID>25</GID>
<name>IN_4</name></connection>
<connection>
<GID>46</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>116 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100.5,-89,-98.5,-89</points>
<connection>
<GID>25</GID>
<name>IN_5</name></connection>
<connection>
<GID>46</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>111 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100.5,-87,-98.5,-87</points>
<connection>
<GID>25</GID>
<name>IN_7</name></connection>
<connection>
<GID>46</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>112 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100.5,-86,-98.5,-86</points>
<connection>
<GID>25</GID>
<name>IN_8</name></connection>
<connection>
<GID>46</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>120 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-100.5,-85,-98.5,-85</points>
<connection>
<GID>25</GID>
<name>IN_9</name></connection>
<connection>
<GID>46</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>422 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-94.5,-96,-94.5,-96</points>
<connection>
<GID>25</GID>
<name>clock</name></connection>
<connection>
<GID>135</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>420 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-98,-77,-98,-76.5</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<intersection>-77 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-98,-77,-94.5,-77</points>
<connection>
<GID>25</GID>
<name>load</name></connection>
<intersection>-98 0</intersection></hsegment></shape></wire>
<wire>
<ID>128 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-93,-45,-93</points>
<connection>
<GID>25</GID>
<name>OUT_1</name></connection>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>-88 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-88,-97.5,-88,-93</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>-93 1</intersection></vsegment></shape></wire>
<wire>
<ID>136 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-84,-45,-84</points>
<connection>
<GID>25</GID>
<name>OUT_10</name></connection>
<connection>
<GID>50</GID>
<name>IN_10</name></connection>
<intersection>-73.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-73.5,-99.5,-73.5,-84</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<intersection>-84 1</intersection></vsegment></shape></wire>
<wire>
<ID>125 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-83,-45,-83</points>
<connection>
<GID>25</GID>
<name>OUT_11</name></connection>
<connection>
<GID>50</GID>
<name>IN_11</name></connection>
<intersection>-73 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-73,-101.5,-73,-83</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>-83 1</intersection></vsegment></shape></wire>
<wire>
<ID>140 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-82,-45,-82</points>
<connection>
<GID>25</GID>
<name>OUT_12</name></connection>
<connection>
<GID>50</GID>
<name>IN_12</name></connection>
<intersection>-66.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-66.5,-95.5,-66.5,-82</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>-82 1</intersection></vsegment></shape></wire>
<wire>
<ID>127 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-81,-45,-81</points>
<connection>
<GID>25</GID>
<name>OUT_13</name></connection>
<connection>
<GID>50</GID>
<name>IN_13</name></connection>
<intersection>-66 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-66,-97.5,-66,-81</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>-81 1</intersection></vsegment></shape></wire>
<wire>
<ID>137 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-80,-45,-80</points>
<connection>
<GID>25</GID>
<name>OUT_14</name></connection>
<connection>
<GID>50</GID>
<name>IN_14</name></connection>
<intersection>-65.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-65.5,-99.5,-65.5,-80</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>-80 1</intersection></vsegment></shape></wire>
<wire>
<ID>300 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-98.5,-123.5,-98.5,-123.5</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<connection>
<GID>88</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>139 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-79,-45,-79</points>
<connection>
<GID>25</GID>
<name>OUT_15</name></connection>
<connection>
<GID>50</GID>
<name>IN_15</name></connection>
<intersection>-65 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-65,-101.5,-65,-79</points>
<connection>
<GID>184</GID>
<name>IN_0</name></connection>
<intersection>-79 1</intersection></vsegment></shape></wire>
<wire>
<ID>130 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-92,-45,-92</points>
<connection>
<GID>25</GID>
<name>OUT_2</name></connection>
<connection>
<GID>50</GID>
<name>IN_2</name></connection>
<intersection>-87.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-87.5,-99.5,-87.5,-92</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>-92 1</intersection></vsegment></shape></wire>
<wire>
<ID>131 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-91,-45,-91</points>
<connection>
<GID>25</GID>
<name>OUT_3</name></connection>
<connection>
<GID>50</GID>
<name>IN_3</name></connection>
<intersection>-87 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-87,-101.5,-87,-91</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>-91 1</intersection></vsegment></shape></wire>
<wire>
<ID>126 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-90,-45,-90</points>
<connection>
<GID>25</GID>
<name>OUT_4</name></connection>
<connection>
<GID>50</GID>
<name>IN_4</name></connection>
<intersection>-81.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-81.5,-95.5,-81.5,-90</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>-90 1</intersection></vsegment></shape></wire>
<wire>
<ID>134 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-89,-45,-89</points>
<connection>
<GID>25</GID>
<name>OUT_5</name></connection>
<connection>
<GID>50</GID>
<name>IN_5</name></connection>
<intersection>-81 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-81,-97.5,-81,-89</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>-89 1</intersection></vsegment></shape></wire>
<wire>
<ID>132 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-87,-45,-87</points>
<connection>
<GID>25</GID>
<name>OUT_7</name></connection>
<connection>
<GID>50</GID>
<name>IN_7</name></connection>
<intersection>-80 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-80,-101.5,-80,-87</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>-87 1</intersection></vsegment></shape></wire>
<wire>
<ID>133 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-86,-45,-86</points>
<connection>
<GID>25</GID>
<name>OUT_8</name></connection>
<connection>
<GID>50</GID>
<name>IN_8</name></connection>
<intersection>-74.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-74.5,-95.5,-74.5,-86</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<intersection>-86 1</intersection></vsegment></shape></wire>
<wire>
<ID>138 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-85,-45,-85</points>
<connection>
<GID>25</GID>
<name>OUT_9</name></connection>
<connection>
<GID>50</GID>
<name>IN_9</name></connection>
<intersection>-74 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-74,-97.5,-74,-85</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>-85 1</intersection></vsegment></shape></wire>
<wire>
<ID>149 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41,-86,-36.5,-86</points>
<connection>
<GID>50</GID>
<name>OUT_8</name></connection>
<connection>
<GID>48</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>302 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-98.5,-121.5,-98.5,-121.5</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<connection>
<GID>27</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>303 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-108.5,-120.5,-98.5,-120.5</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<connection>
<GID>27</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>157 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-114.5,-49,-114.5</points>
<connection>
<GID>52</GID>
<name>IN_9</name></connection>
<connection>
<GID>27</GID>
<name>OUT_9</name></connection>
<intersection>-74 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-74,-127,-74,-114.5</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<intersection>-114.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>310 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-98.5,-113.5,-98.5,-113.5</points>
<connection>
<GID>27</GID>
<name>IN_10</name></connection>
<connection>
<GID>98</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>311 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-108.5,-112.5,-98.5,-112.5</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<connection>
<GID>27</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>167 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-121.5,-49,-121.5</points>
<connection>
<GID>52</GID>
<name>IN_2</name></connection>
<connection>
<GID>27</GID>
<name>OUT_2</name></connection>
<intersection>-87.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-87.5,-129,-87.5,-121.5</points>
<connection>
<GID>189</GID>
<name>IN_0</name></connection>
<intersection>-121.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>312 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-98.5,-111.5,-98.5,-111.5</points>
<connection>
<GID>27</GID>
<name>IN_12</name></connection>
<connection>
<GID>100</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>313 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-108.5,-110.5,-98.5,-110.5</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<connection>
<GID>27</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>161 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-122.5,-49,-122.5</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<connection>
<GID>27</GID>
<name>OUT_1</name></connection>
<intersection>-88 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-88,-127,-88,-122.5</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>-122.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>314 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-98.5,-109.5,-98.5,-109.5</points>
<connection>
<GID>27</GID>
<name>IN_14</name></connection>
<connection>
<GID>102</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>315 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-108.5,-108.5,-98.5,-108.5</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<connection>
<GID>27</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>159 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-119.5,-49,-119.5</points>
<connection>
<GID>52</GID>
<name>IN_4</name></connection>
<connection>
<GID>27</GID>
<name>OUT_4</name></connection>
<intersection>-81.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-81.5,-125,-81.5,-119.5</points>
<connection>
<GID>191</GID>
<name>IN_0</name></connection>
<intersection>-119.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>304 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-98.5,-119.5,-98.5,-119.5</points>
<connection>
<GID>27</GID>
<name>IN_4</name></connection>
<connection>
<GID>92</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>305 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-108.5,-118.5,-98.5,-118.5</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<connection>
<GID>27</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>306 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-98.5,-117.5,-98.5,-117.5</points>
<connection>
<GID>27</GID>
<name>IN_6</name></connection>
<connection>
<GID>94</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>307 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-108.5,-116.5,-98.5,-116.5</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<connection>
<GID>27</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>147 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41,-90,-36.5,-90</points>
<connection>
<GID>50</GID>
<name>OUT_4</name></connection>
<connection>
<GID>48</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>308 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-98.5,-115.5,-98.5,-115.5</points>
<connection>
<GID>27</GID>
<name>IN_8</name></connection>
<connection>
<GID>96</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>309 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-108.5,-114.5,-98.5,-114.5</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<connection>
<GID>27</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>426 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-92.5,-125.5,-92.5,-125.5</points>
<connection>
<GID>27</GID>
<name>clear</name></connection>
<connection>
<GID>143</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>425 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-94.5,-125.5,-94.5,-125.5</points>
<connection>
<GID>27</GID>
<name>clock</name></connection>
<connection>
<GID>141</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>424 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-89.5,-106.5,-89.5,-104.5</points>
<connection>
<GID>139</GID>
<name>IN_0</name></connection>
<intersection>-106.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-93.5,-106.5,-89.5,-106.5</points>
<connection>
<GID>27</GID>
<name>count_enable</name></connection>
<intersection>-89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>164 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-123.5,-49,-123.5</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>-88.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-88.5,-125,-88.5,-123.5</points>
<connection>
<GID>186</GID>
<name>IN_0</name></connection>
<intersection>-123.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1033 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-51,-27.5,-42,-27.5</points>
<connection>
<GID>107</GID>
<name>OUT_13</name></connection>
<connection>
<GID>109</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>318 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-59.5,-38.5,-55,-38.5</points>
<connection>
<GID>105</GID>
<name>IN_2</name></connection>
<connection>
<GID>107</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>165 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-113.5,-49,-113.5</points>
<connection>
<GID>52</GID>
<name>IN_10</name></connection>
<connection>
<GID>27</GID>
<name>OUT_10</name></connection>
<intersection>-73.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-73.5,-129,-73.5,-113.5</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<intersection>-113.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>166 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-112.5,-49,-112.5</points>
<connection>
<GID>52</GID>
<name>IN_11</name></connection>
<connection>
<GID>27</GID>
<name>OUT_11</name></connection>
<intersection>-73 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-73,-131,-73,-112.5</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>-112.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>158 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-111.5,-49,-111.5</points>
<connection>
<GID>52</GID>
<name>IN_12</name></connection>
<connection>
<GID>27</GID>
<name>OUT_12</name></connection>
<intersection>-66.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-66.5,-125,-66.5,-111.5</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<intersection>-111.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1040 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-59.5,-26.5,-55,-26.5</points>
<connection>
<GID>107</GID>
<name>IN_14</name></connection>
<connection>
<GID>105</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>172 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-110.5,-49,-110.5</points>
<connection>
<GID>52</GID>
<name>IN_13</name></connection>
<connection>
<GID>27</GID>
<name>OUT_13</name></connection>
<intersection>-66 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-66,-127,-66,-110.5</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<intersection>-110.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>163 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-109.5,-49,-109.5</points>
<connection>
<GID>52</GID>
<name>IN_14</name></connection>
<connection>
<GID>27</GID>
<name>OUT_14</name></connection>
<intersection>-65.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-65.5,-129,-65.5,-109.5</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<intersection>-109.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>170 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-108.5,-49,-108.5</points>
<connection>
<GID>52</GID>
<name>IN_15</name></connection>
<connection>
<GID>27</GID>
<name>OUT_15</name></connection>
<intersection>-65 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-65,-131,-65,-108.5</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>-108.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>160 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-120.5,-49,-120.5</points>
<connection>
<GID>52</GID>
<name>IN_3</name></connection>
<connection>
<GID>27</GID>
<name>OUT_3</name></connection>
<intersection>-87 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-87,-131,-87,-120.5</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<intersection>-120.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>171 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-117.5,-49,-117.5</points>
<connection>
<GID>52</GID>
<name>IN_6</name></connection>
<connection>
<GID>27</GID>
<name>OUT_6</name></connection>
<intersection>-80.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-80.5,-129,-80.5,-117.5</points>
<connection>
<GID>193</GID>
<name>IN_0</name></connection>
<intersection>-117.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>162 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-116.5,-49,-116.5</points>
<connection>
<GID>52</GID>
<name>IN_7</name></connection>
<connection>
<GID>27</GID>
<name>OUT_7</name></connection>
<intersection>-80 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-80,-131,-80,-116.5</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>-116.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>168 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-88.5,-115.5,-49,-115.5</points>
<connection>
<GID>52</GID>
<name>IN_8</name></connection>
<connection>
<GID>27</GID>
<name>OUT_8</name></connection>
<intersection>-74.5 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-74.5,-125,-74.5,-115.5</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>-115.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>190 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-104.5,-154,-99,-154</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<connection>
<GID>58</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>191 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-104.5,-153,-99,-153</points>
<connection>
<GID>29</GID>
<name>IN_1</name></connection>
<connection>
<GID>58</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>197 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-104.5,-144,-99,-144</points>
<connection>
<GID>29</GID>
<name>IN_10</name></connection>
<connection>
<GID>58</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>200 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-104.5,-143,-99,-143</points>
<connection>
<GID>29</GID>
<name>IN_11</name></connection>
<connection>
<GID>58</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>204 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-104.5,-142,-99,-142</points>
<connection>
<GID>29</GID>
<name>IN_12</name></connection>
<connection>
<GID>58</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>199 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-104.5,-141,-99,-141</points>
<connection>
<GID>29</GID>
<name>IN_13</name></connection>
<connection>
<GID>58</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>201 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-104.5,-139,-99,-139</points>
<connection>
<GID>29</GID>
<name>IN_15</name></connection>
<connection>
<GID>58</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>189 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-104.5,-152,-99,-152</points>
<connection>
<GID>29</GID>
<name>IN_2</name></connection>
<connection>
<GID>58</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>192 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-104.5,-151,-99,-151</points>
<connection>
<GID>29</GID>
<name>IN_3</name></connection>
<connection>
<GID>58</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>194 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-104.5,-150,-99,-150</points>
<connection>
<GID>29</GID>
<name>IN_4</name></connection>
<connection>
<GID>58</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>196 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-104.5,-149,-99,-149</points>
<connection>
<GID>29</GID>
<name>IN_5</name></connection>
<connection>
<GID>58</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>195 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-104.5,-148,-99,-148</points>
<connection>
<GID>29</GID>
<name>IN_6</name></connection>
<connection>
<GID>58</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>346 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-51,-39.5,-42,-39.5</points>
<connection>
<GID>109</GID>
<name>IN_1</name></connection>
<connection>
<GID>107</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>193 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-104.5,-147,-99,-147</points>
<connection>
<GID>29</GID>
<name>IN_7</name></connection>
<connection>
<GID>58</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>198 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-104.5,-146,-99,-146</points>
<connection>
<GID>29</GID>
<name>IN_8</name></connection>
<connection>
<GID>58</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>202 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-104.5,-145,-99,-145</points>
<connection>
<GID>29</GID>
<name>IN_9</name></connection>
<connection>
<GID>58</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>427 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-98,-137,-95,-137</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<connection>
<GID>29</GID>
<name>load</name></connection></hsegment></shape></wire>
<wire>
<ID>219 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89,-154,-46,-154</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>-89 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-89,-155.5,-89,-154</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<intersection>-154 1</intersection></vsegment></shape></wire>
<wire>
<ID>209 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89,-153,-46,-153</points>
<connection>
<GID>29</GID>
<name>OUT_1</name></connection>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<intersection>-88.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-88.5,-157.5,-88.5,-153</points>
<connection>
<GID>204</GID>
<name>IN_0</name></connection>
<intersection>-153 1</intersection></vsegment></shape></wire>
<wire>
<ID>218 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89,-144,-46,-144</points>
<connection>
<GID>29</GID>
<name>OUT_10</name></connection>
<connection>
<GID>62</GID>
<name>IN_10</name></connection>
<intersection>-68 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-68,-159.5,-68,-144</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>-144 1</intersection></vsegment></shape></wire>
<wire>
<ID>550 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41,-79,-36.5,-79</points>
<connection>
<GID>48</GID>
<name>IN_15</name></connection>
<connection>
<GID>50</GID>
<name>OUT_15</name></connection></hsegment></shape></wire>
<wire>
<ID>220 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89,-143,-46,-143</points>
<connection>
<GID>29</GID>
<name>OUT_11</name></connection>
<connection>
<GID>62</GID>
<name>IN_11</name></connection>
<intersection>-67.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-67.5,-161.5,-67.5,-143</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<intersection>-143 1</intersection></vsegment></shape></wire>
<wire>
<ID>205 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89,-142,-46,-142</points>
<connection>
<GID>29</GID>
<name>OUT_12</name></connection>
<connection>
<GID>62</GID>
<name>IN_12</name></connection>
<intersection>-62 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-62,-155.5,-62,-142</points>
<connection>
<GID>215</GID>
<name>IN_0</name></connection>
<intersection>-142 1</intersection></vsegment></shape></wire>
<wire>
<ID>207 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89,-141,-46,-141</points>
<connection>
<GID>29</GID>
<name>OUT_13</name></connection>
<connection>
<GID>62</GID>
<name>IN_13</name></connection>
<intersection>-61.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-61.5,-157.5,-61.5,-141</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<intersection>-141 1</intersection></vsegment></shape></wire>
<wire>
<ID>206 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89,-140,-46,-140</points>
<connection>
<GID>62</GID>
<name>IN_14</name></connection>
<connection>
<GID>29</GID>
<name>OUT_14</name></connection>
<intersection>-60.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-60.5,-159.5,-60.5,-140</points>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<intersection>-140 1</intersection></vsegment></shape></wire>
<wire>
<ID>208 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89,-139,-46,-139</points>
<connection>
<GID>29</GID>
<name>OUT_15</name></connection>
<connection>
<GID>62</GID>
<name>IN_15</name></connection>
<intersection>-60 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-60,-161.5,-60,-139</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<intersection>-139 1</intersection></vsegment></shape></wire>
<wire>
<ID>210 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89,-152,-46,-152</points>
<connection>
<GID>29</GID>
<name>OUT_2</name></connection>
<connection>
<GID>62</GID>
<name>IN_2</name></connection>
<intersection>-88 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-88,-159.5,-88,-152</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<intersection>-152 1</intersection></vsegment></shape></wire>
<wire>
<ID>212 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89,-150,-46,-150</points>
<connection>
<GID>29</GID>
<name>OUT_4</name></connection>
<connection>
<GID>62</GID>
<name>IN_4</name></connection>
<intersection>-83 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-83,-155.5,-83,-150</points>
<connection>
<GID>207</GID>
<name>IN_0</name></connection>
<intersection>-150 1</intersection></vsegment></shape></wire>
<wire>
<ID>214 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89,-148,-46,-148</points>
<connection>
<GID>29</GID>
<name>OUT_6</name></connection>
<connection>
<GID>62</GID>
<name>IN_6</name></connection>
<intersection>-82 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-82,-159.5,-82,-148</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<intersection>-148 1</intersection></vsegment></shape></wire>
<wire>
<ID>215 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89,-147,-46,-147</points>
<connection>
<GID>29</GID>
<name>OUT_7</name></connection>
<connection>
<GID>62</GID>
<name>IN_7</name></connection>
<intersection>-81.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-81.5,-161.5,-81.5,-147</points>
<connection>
<GID>210</GID>
<name>IN_0</name></connection>
<intersection>-147 1</intersection></vsegment></shape></wire>
<wire>
<ID>216 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-89,-146,-46,-146</points>
<connection>
<GID>29</GID>
<name>OUT_8</name></connection>
<connection>
<GID>62</GID>
<name>IN_8</name></connection>
<intersection>-69 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-69,-155.5,-69,-146</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<intersection>-146 1</intersection></vsegment></shape></wire>
<wire>
<ID>238 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-105.5,-180,-99.5,-180</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<connection>
<GID>66</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>248 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-105.5,-171,-99.5,-171</points>
<connection>
<GID>31</GID>
<name>IN_10</name></connection>
<connection>
<GID>66</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>242 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-105.5,-167,-99.5,-167</points>
<connection>
<GID>31</GID>
<name>IN_14</name></connection>
<connection>
<GID>66</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>240 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-105.5,-179,-99.5,-179</points>
<connection>
<GID>31</GID>
<name>IN_2</name></connection>
<connection>
<GID>66</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>246 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-105.5,-175,-99.5,-175</points>
<connection>
<GID>31</GID>
<name>IN_6</name></connection>
<connection>
<GID>66</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>250 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-105.5,-174,-99.5,-174</points>
<connection>
<GID>31</GID>
<name>IN_7</name></connection>
<connection>
<GID>66</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>252 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-105.5,-173,-99.5,-173</points>
<connection>
<GID>31</GID>
<name>IN_8</name></connection>
<connection>
<GID>66</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>244 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-105.5,-172,-99.5,-172</points>
<connection>
<GID>31</GID>
<name>IN_9</name></connection>
<connection>
<GID>66</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>432 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-95.5,-183,-95.5,-183</points>
<connection>
<GID>31</GID>
<name>clock</name></connection>
<connection>
<GID>155</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>430 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-97.5,-164,-95.5,-164</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<connection>
<GID>31</GID>
<name>load</name></connection></hsegment></shape></wire>
<wire>
<ID>1061 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-87,-23.5,-84,-23.5</points>
<connection>
<GID>539</GID>
<name>OUT_0</name></connection>
<intersection>-84 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-84,-28.5,-84,-23.5</points>
<connection>
<GID>38</GID>
<name>IN_12</name></connection>
<connection>
<GID>38</GID>
<name>IN_13</name></connection>
<connection>
<GID>38</GID>
<name>IN_14</name></connection>
<connection>
<GID>38</GID>
<name>IN_15</name></connection>
<intersection>-23.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>82 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-80.5,-65.5,-77.5,-65.5</points>
<connection>
<GID>42</GID>
<name>Bus_in_0</name></connection>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>83 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-80.5,-64.5,-77.5,-64.5</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<connection>
<GID>44</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>101 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-80.5,-55.5,-77.5,-55.5</points>
<connection>
<GID>42</GID>
<name>IN_10</name></connection>
<connection>
<GID>44</GID>
<name>OUT_10</name></connection></hsegment></shape></wire>
<wire>
<ID>103 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-80.5,-54.5,-77.5,-54.5</points>
<connection>
<GID>42</GID>
<name>IN_11</name></connection>
<connection>
<GID>44</GID>
<name>OUT_11</name></connection></hsegment></shape></wire>
<wire>
<ID>108 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-80.5,-63.5,-77.5,-63.5</points>
<connection>
<GID>42</GID>
<name>IN_2</name></connection>
<connection>
<GID>44</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>100 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-80.5,-62.5,-77.5,-62.5</points>
<connection>
<GID>42</GID>
<name>IN_3</name></connection>
<connection>
<GID>44</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>105 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-80.5,-61.5,-77.5,-61.5</points>
<connection>
<GID>42</GID>
<name>IN_4</name></connection>
<connection>
<GID>44</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>102 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-80.5,-60.5,-77.5,-60.5</points>
<connection>
<GID>42</GID>
<name>IN_5</name></connection>
<connection>
<GID>44</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>106 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-80.5,-59.5,-77.5,-59.5</points>
<connection>
<GID>42</GID>
<name>IN_6</name></connection>
<connection>
<GID>44</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>98 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-80.5,-58.5,-77.5,-58.5</points>
<connection>
<GID>42</GID>
<name>IN_7</name></connection>
<connection>
<GID>44</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>99 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-80.5,-57.5,-77.5,-57.5</points>
<connection>
<GID>42</GID>
<name>IN_8</name></connection>
<connection>
<GID>44</GID>
<name>OUT_8</name></connection></hsegment></shape></wire>
<wire>
<ID>107 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-80.5,-56.5,-77.5,-56.5</points>
<connection>
<GID>42</GID>
<name>IN_9</name></connection>
<connection>
<GID>44</GID>
<name>OUT_9</name></connection></hsegment></shape></wire>
<wire>
<ID>434 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-79,-49,-79,-48.5</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>-49 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-82.5,-49,-79,-49</points>
<connection>
<GID>44</GID>
<name>ENABLE_0</name></connection>
<intersection>-79 0</intersection></hsegment></shape></wire>
<wire>
<ID>143 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41,-94,-36.5,-94</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<connection>
<GID>48</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>144 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41,-93,-36.5,-93</points>
<connection>
<GID>50</GID>
<name>OUT_1</name></connection>
<connection>
<GID>48</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>152 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41,-84,-36.5,-84</points>
<connection>
<GID>50</GID>
<name>OUT_10</name></connection>
<connection>
<GID>48</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>156 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41,-83,-36.5,-83</points>
<connection>
<GID>50</GID>
<name>OUT_11</name></connection>
<connection>
<GID>48</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>543 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41,-82,-36.5,-82</points>
<connection>
<GID>50</GID>
<name>OUT_12</name></connection>
<connection>
<GID>48</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>548 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41,-80,-36.5,-80</points>
<connection>
<GID>50</GID>
<name>OUT_14</name></connection>
<connection>
<GID>48</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>146 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41,-92,-36.5,-92</points>
<connection>
<GID>50</GID>
<name>OUT_2</name></connection>
<connection>
<GID>48</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>145 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41,-91,-36.5,-91</points>
<connection>
<GID>50</GID>
<name>OUT_3</name></connection>
<connection>
<GID>48</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>141 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41,-89,-36.5,-89</points>
<connection>
<GID>50</GID>
<name>OUT_5</name></connection>
<connection>
<GID>48</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>142 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41,-88,-36.5,-88</points>
<connection>
<GID>50</GID>
<name>OUT_6</name></connection>
<connection>
<GID>48</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>154 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41,-87,-36.5,-87</points>
<connection>
<GID>50</GID>
<name>OUT_7</name></connection>
<connection>
<GID>48</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1039 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-59.5,-27.5,-55,-27.5</points>
<connection>
<GID>105</GID>
<name>IN_13</name></connection>
<connection>
<GID>107</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>316 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-59.5,-40.5,-55,-40.5</points>
<connection>
<GID>105</GID>
<name>Bus_in_0</name></connection>
<connection>
<GID>107</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>155 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41,-85,-36.5,-85</points>
<connection>
<GID>50</GID>
<name>OUT_9</name></connection>
<connection>
<GID>48</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>435 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-77.5,-43,-77.5</points>
<connection>
<GID>50</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>161</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>436 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-47,-107,-47,-107</points>
<connection>
<GID>52</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>163</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>182 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-45,-123.5,-36.5,-123.5</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<connection>
<GID>56</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>177 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-45,-122.5,-36.5,-122.5</points>
<connection>
<GID>52</GID>
<name>OUT_1</name></connection>
<connection>
<GID>56</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>176 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-45,-113.5,-36.5,-113.5</points>
<connection>
<GID>52</GID>
<name>OUT_10</name></connection>
<connection>
<GID>56</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>174 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-45,-112.5,-36.5,-112.5</points>
<connection>
<GID>52</GID>
<name>OUT_11</name></connection>
<connection>
<GID>56</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>178 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-45,-111.5,-36.5,-111.5</points>
<connection>
<GID>52</GID>
<name>OUT_12</name></connection>
<connection>
<GID>56</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>180 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-45,-110.5,-36.5,-110.5</points>
<connection>
<GID>52</GID>
<name>OUT_13</name></connection>
<connection>
<GID>56</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>181 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-45,-109.5,-36.5,-109.5</points>
<connection>
<GID>52</GID>
<name>OUT_14</name></connection>
<connection>
<GID>56</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>183 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-45,-108.5,-36.5,-108.5</points>
<connection>
<GID>52</GID>
<name>OUT_15</name></connection>
<connection>
<GID>56</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>173 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-45,-121.5,-36.5,-121.5</points>
<connection>
<GID>52</GID>
<name>OUT_2</name></connection>
<connection>
<GID>56</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>188 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-45,-120.5,-36.5,-120.5</points>
<connection>
<GID>52</GID>
<name>OUT_3</name></connection>
<connection>
<GID>56</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>186 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-45,-119.5,-36.5,-119.5</points>
<connection>
<GID>52</GID>
<name>OUT_4</name></connection>
<connection>
<GID>56</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>179 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-45,-117.5,-36.5,-117.5</points>
<connection>
<GID>52</GID>
<name>OUT_6</name></connection>
<connection>
<GID>56</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>185 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-45,-116.5,-36.5,-116.5</points>
<connection>
<GID>52</GID>
<name>OUT_7</name></connection>
<connection>
<GID>56</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>175 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-45,-115.5,-36.5,-115.5</points>
<connection>
<GID>52</GID>
<name>OUT_8</name></connection>
<connection>
<GID>56</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>187 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-45,-114.5,-36.5,-114.5</points>
<connection>
<GID>52</GID>
<name>OUT_9</name></connection>
<connection>
<GID>56</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>228 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-42,-154,-36.5,-154</points>
<connection>
<GID>60</GID>
<name>Bus_in_0</name></connection>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>232 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-42,-153,-36.5,-153</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<connection>
<GID>62</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>224 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-42,-143,-36.5,-143</points>
<connection>
<GID>60</GID>
<name>IN_11</name></connection>
<connection>
<GID>62</GID>
<name>OUT_11</name></connection></hsegment></shape></wire>
<wire>
<ID>226 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-42,-141,-36.5,-141</points>
<connection>
<GID>60</GID>
<name>IN_13</name></connection>
<connection>
<GID>62</GID>
<name>OUT_13</name></connection></hsegment></shape></wire>
<wire>
<ID>236 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-42,-140,-36.5,-140</points>
<connection>
<GID>60</GID>
<name>IN_14</name></connection>
<connection>
<GID>62</GID>
<name>OUT_14</name></connection></hsegment></shape></wire>
<wire>
<ID>222 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-42,-151,-36.5,-151</points>
<connection>
<GID>60</GID>
<name>IN_3</name></connection>
<connection>
<GID>62</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>229 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-42,-149,-36.5,-149</points>
<connection>
<GID>60</GID>
<name>IN_5</name></connection>
<connection>
<GID>62</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>234 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-42,-147,-36.5,-147</points>
<connection>
<GID>60</GID>
<name>IN_7</name></connection>
<connection>
<GID>62</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>230 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-42,-146,-36.5,-146</points>
<connection>
<GID>60</GID>
<name>IN_8</name></connection>
<connection>
<GID>62</GID>
<name>OUT_8</name></connection></hsegment></shape></wire>
<wire>
<ID>437 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-44,-137.5,-44,-137.5</points>
<connection>
<GID>62</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>165</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>324 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-59.5,-30.5,-55,-30.5</points>
<connection>
<GID>105</GID>
<name>IN_10</name></connection>
<connection>
<GID>107</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>1038 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-59.5,-28.5,-55,-28.5</points>
<connection>
<GID>107</GID>
<name>IN_12</name></connection>
<connection>
<GID>105</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>1044 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-59.5,-25.5,-55,-25.5</points>
<connection>
<GID>105</GID>
<name>IN_15</name></connection>
<connection>
<GID>107</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>319 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-59.5,-37.5,-55,-37.5</points>
<connection>
<GID>105</GID>
<name>IN_3</name></connection>
<connection>
<GID>107</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>320 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-59.5,-36.5,-55,-36.5</points>
<connection>
<GID>105</GID>
<name>IN_4</name></connection>
<connection>
<GID>107</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>325 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-59.5,-35.5,-55,-35.5</points>
<connection>
<GID>105</GID>
<name>IN_5</name></connection>
<connection>
<GID>107</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>329 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-59.5,-34.5,-55,-34.5</points>
<connection>
<GID>105</GID>
<name>IN_6</name></connection>
<connection>
<GID>107</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>327 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-59.5,-33.5,-55,-33.5</points>
<connection>
<GID>105</GID>
<name>IN_7</name></connection>
<connection>
<GID>107</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>330 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-59.5,-32.5,-55,-32.5</points>
<connection>
<GID>105</GID>
<name>IN_8</name></connection>
<connection>
<GID>107</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>326 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-59.5,-31.5,-55,-31.5</points>
<connection>
<GID>105</GID>
<name>IN_9</name></connection>
<connection>
<GID>107</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>433 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-53,-24,-53,-24</points>
<connection>
<GID>107</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>157</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>337 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-51,-40.5,-42,-40.5</points>
<connection>
<GID>109</GID>
<name>Bus_in_0</name></connection>
<connection>
<GID>107</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>340 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-51,-30.5,-42,-30.5</points>
<connection>
<GID>109</GID>
<name>IN_10</name></connection>
<connection>
<GID>107</GID>
<name>OUT_10</name></connection></hsegment></shape></wire>
<wire>
<ID>342 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-51,-29.5,-42,-29.5</points>
<connection>
<GID>109</GID>
<name>IN_11</name></connection>
<connection>
<GID>107</GID>
<name>OUT_11</name></connection></hsegment></shape></wire>
<wire>
<ID>1027 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-51,-28.5,-42,-28.5</points>
<connection>
<GID>109</GID>
<name>IN_12</name></connection>
<connection>
<GID>107</GID>
<name>OUT_12</name></connection></hsegment></shape></wire>
<wire>
<ID>1036 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-51,-26.5,-42,-26.5</points>
<connection>
<GID>109</GID>
<name>IN_14</name></connection>
<connection>
<GID>107</GID>
<name>OUT_14</name></connection></hsegment></shape></wire>
<wire>
<ID>1037 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-51,-25.5,-42,-25.5</points>
<connection>
<GID>107</GID>
<name>OUT_15</name></connection>
<connection>
<GID>109</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>334 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-51,-38.5,-42,-38.5</points>
<connection>
<GID>109</GID>
<name>IN_2</name></connection>
<connection>
<GID>107</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>335 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-51,-37.5,-42,-37.5</points>
<connection>
<GID>109</GID>
<name>IN_3</name></connection>
<connection>
<GID>107</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>338 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-51,-36.5,-42,-36.5</points>
<connection>
<GID>109</GID>
<name>IN_4</name></connection>
<connection>
<GID>107</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>332 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-51,-35.5,-42,-35.5</points>
<connection>
<GID>109</GID>
<name>IN_5</name></connection>
<connection>
<GID>107</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>336 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-51,-34.5,-42,-34.5</points>
<connection>
<GID>109</GID>
<name>IN_6</name></connection>
<connection>
<GID>107</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>339 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-51,-33.5,-42,-33.5</points>
<connection>
<GID>109</GID>
<name>IN_7</name></connection>
<connection>
<GID>107</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>347 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-51,-32.5,-42,-32.5</points>
<connection>
<GID>109</GID>
<name>IN_8</name></connection>
<connection>
<GID>107</GID>
<name>OUT_8</name></connection></hsegment></shape></wire>
<wire>
<ID>341 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-51,-31.5,-42,-31.5</points>
<connection>
<GID>109</GID>
<name>IN_9</name></connection>
<connection>
<GID>107</GID>
<name>OUT_9</name></connection></hsegment></shape></wire>
<wire>
<ID>410 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-22,21,-22</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<connection>
<GID>111</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>408 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-12,21,-12</points>
<connection>
<GID>113</GID>
<name>IN_10</name></connection>
<connection>
<GID>111</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>396 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-11,21,-11</points>
<connection>
<GID>113</GID>
<name>IN_11</name></connection>
<connection>
<GID>111</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>402 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-9,21,-9</points>
<connection>
<GID>113</GID>
<name>IN_13</name></connection>
<connection>
<GID>111</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>400 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-20,21,-20</points>
<connection>
<GID>113</GID>
<name>IN_2</name></connection>
<connection>
<GID>111</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>398 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-18,21,-18</points>
<connection>
<GID>113</GID>
<name>IN_4</name></connection>
<connection>
<GID>111</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>406 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-15,21,-15</points>
<connection>
<GID>113</GID>
<name>IN_7</name></connection>
<connection>
<GID>111</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>404 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-14,21,-14</points>
<connection>
<GID>113</GID>
<name>IN_8</name></connection>
<connection>
<GID>111</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>412 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-25,25,-24</points>
<connection>
<GID>113</GID>
<name>clock</name></connection>
<connection>
<GID>115</GID>
<name>IN_0</name></connection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>39.0819,-2.02822,225.425,-94.5326</PageViewport>
<gate>
<ID>77</ID>
<type>DE_TO</type>
<position>67,-55</position>
<input>
<ID>IN_0</ID>440 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add11</lparam></gate>
<gate>
<ID>13</ID>
<type>DE_TO</type>
<position>67,-19</position>
<input>
<ID>IN_0</ID>71 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add2</lparam></gate>
<gate>
<ID>69</ID>
<type>DE_TO</type>
<position>67,-53</position>
<input>
<ID>IN_0</ID>439 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add10</lparam></gate>
<gate>
<ID>5</ID>
<type>AE_FULLADDER_4BIT</type>
<position>61,-18</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>79 </input>
<input>
<ID>IN_2</ID>80 </input>
<input>
<ID>IN_3</ID>285 </input>
<input>
<ID>IN_B_0</ID>77 </input>
<input>
<ID>IN_B_1</ID>74 </input>
<input>
<ID>IN_B_2</ID>75 </input>
<input>
<ID>IN_B_3</ID>76 </input>
<output>
<ID>OUT_0</ID>69 </output>
<output>
<ID>OUT_1</ID>70 </output>
<output>
<ID>OUT_2</ID>71 </output>
<output>
<ID>OUT_3</ID>72 </output>
<input>
<ID>carry_in</ID>465 </input>
<output>
<ID>carry_out</ID>461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>33</ID>
<type>DA_FROM</type>
<position>55,-17.5</position>
<input>
<ID>IN_0</ID>76 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr3</lparam></gate>
<gate>
<ID>735</ID>
<type>DA_FROM</type>
<position>243.5,-186</position>
<input>
<ID>IN_0</ID>979 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr15</lparam></gate>
<gate>
<ID>73</ID>
<type>DE_TO</type>
<position>67,-49</position>
<input>
<ID>IN_0</ID>298 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add8</lparam></gate>
<gate>
<ID>9</ID>
<type>DE_TO</type>
<position>67,-15</position>
<input>
<ID>IN_0</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add0</lparam></gate>
<gate>
<ID>711</ID>
<type>DA_FROM</type>
<position>88.5,-186</position>
<input>
<ID>IN_0</ID>955 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr12</lparam></gate>
<gate>
<ID>75</ID>
<type>DE_TO</type>
<position>67,-51</position>
<input>
<ID>IN_0</ID>299 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add9</lparam></gate>
<gate>
<ID>11</ID>
<type>DE_TO</type>
<position>67,-17</position>
<input>
<ID>IN_0</ID>70 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add1</lparam></gate>
<gate>
<ID>35</ID>
<type>DA_FROM</type>
<position>55,-11.5</position>
<input>
<ID>IN_0</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr0</lparam></gate>
<gate>
<ID>24</ID>
<type>DA_FROM</type>
<position>55,-15.5</position>
<input>
<ID>IN_0</ID>75 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr2</lparam></gate>
<gate>
<ID>80</ID>
<type>DA_FROM</type>
<position>55,-56</position>
<input>
<ID>IN_0</ID>446 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac9</lparam></gate>
<gate>
<ID>511</ID>
<type>AA_AND2</type>
<position>248.5,-165.5</position>
<input>
<ID>IN_0</ID>762 </input>
<input>
<ID>IN_1</ID>763 </input>
<output>
<ID>OUT</ID>775 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>DE_TO</type>
<position>67,-21</position>
<input>
<ID>IN_0</ID>72 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add3</lparam></gate>
<gate>
<ID>84</ID>
<type>AE_FULLADDER_4BIT</type>
<position>61,-69</position>
<input>
<ID>IN_0</ID>457 </input>
<input>
<ID>IN_1</ID>458 </input>
<input>
<ID>IN_2</ID>459 </input>
<input>
<ID>IN_3</ID>460 </input>
<input>
<ID>IN_B_0</ID>456 </input>
<input>
<ID>IN_B_1</ID>453 </input>
<input>
<ID>IN_B_2</ID>454 </input>
<input>
<ID>IN_B_3</ID>455 </input>
<output>
<ID>OUT_0</ID>449 </output>
<output>
<ID>OUT_1</ID>450 </output>
<output>
<ID>OUT_2</ID>451 </output>
<output>
<ID>OUT_3</ID>452 </output>
<input>
<ID>carry_in</ID>463 </input>
<output>
<ID>carry_out</ID>464 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>499</ID>
<type>AE_SMALL_INVERTER</type>
<position>192,-166.5</position>
<input>
<ID>IN_0</ID>944 </input>
<output>
<ID>OUT_0</ID>739 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>20</ID>
<type>DA_FROM</type>
<position>55,-13.5</position>
<input>
<ID>IN_0</ID>74 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr1</lparam></gate>
<gate>
<ID>723</ID>
<type>DA_FROM</type>
<position>140,-206</position>
<input>
<ID>IN_0</ID>967 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr13</lparam></gate>
<gate>
<ID>37</ID>
<type>DA_FROM</type>
<position>55,-20</position>
<input>
<ID>IN_0</ID>78 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac0</lparam></gate>
<gate>
<ID>743</ID>
<type>DE_TO</type>
<position>229,-69.5</position>
<input>
<ID>IN_0</ID>987 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN2</lparam></gate>
<gate>
<ID>41</ID>
<type>DA_FROM</type>
<position>55,-22</position>
<input>
<ID>IN_0</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac1</lparam></gate>
<gate>
<ID>43</ID>
<type>DA_FROM</type>
<position>55,-24</position>
<input>
<ID>IN_0</ID>80 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac2</lparam></gate>
<gate>
<ID>731</ID>
<type>DA_FROM</type>
<position>192,-206</position>
<input>
<ID>IN_0</ID>975 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr14</lparam></gate>
<gate>
<ID>45</ID>
<type>DA_FROM</type>
<position>55,-26</position>
<input>
<ID>IN_0</ID>285 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac3</lparam></gate>
<gate>
<ID>47</ID>
<type>DE_TO</type>
<position>67,-36</position>
<input>
<ID>IN_0</ID>288 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add6</lparam></gate>
<gate>
<ID>751</ID>
<type>DE_TO</type>
<position>228.5,-160</position>
<input>
<ID>IN_0</ID>995 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN10</lparam></gate>
<gate>
<ID>49</ID>
<type>AE_FULLADDER_4BIT</type>
<position>61,-35</position>
<input>
<ID>IN_0</ID>294 </input>
<input>
<ID>IN_1</ID>295 </input>
<input>
<ID>IN_2</ID>296 </input>
<input>
<ID>IN_3</ID>297 </input>
<input>
<ID>IN_B_0</ID>293 </input>
<input>
<ID>IN_B_1</ID>290 </input>
<input>
<ID>IN_B_2</ID>291 </input>
<input>
<ID>IN_B_3</ID>292 </input>
<output>
<ID>OUT_0</ID>286 </output>
<output>
<ID>OUT_1</ID>287 </output>
<output>
<ID>OUT_2</ID>288 </output>
<output>
<ID>OUT_3</ID>289 </output>
<input>
<ID>carry_in</ID>461 </input>
<output>
<ID>carry_out</ID>462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>51</ID>
<type>DA_FROM</type>
<position>55,-34.5</position>
<input>
<ID>IN_0</ID>292 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr7</lparam></gate>
<gate>
<ID>739</ID>
<type>DA_FROM</type>
<position>243.5,-206</position>
<input>
<ID>IN_0</ID>983 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr15</lparam></gate>
<gate>
<ID>53</ID>
<type>DE_TO</type>
<position>67,-32</position>
<input>
<ID>IN_0</ID>286 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add4</lparam></gate>
<gate>
<ID>477</ID>
<type>AE_SMALL_INVERTER</type>
<position>140,-166.5</position>
<input>
<ID>IN_0</ID>936 </input>
<output>
<ID>OUT_0</ID>715 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>118</ID>
<type>DA_FROM</type>
<position>55,-77</position>
<input>
<ID>IN_0</ID>460 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac15</lparam></gate>
<gate>
<ID>748</ID>
<type>DE_TO</type>
<position>280.5,-115</position>
<input>
<ID>IN_0</ID>992 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN7</lparam></gate>
<gate>
<ID>54</ID>
<type>DA_FROM</type>
<position>55,-28.5</position>
<input>
<ID>IN_0</ID>293 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr4</lparam></gate>
<gate>
<ID>55</ID>
<type>DE_TO</type>
<position>67,-34</position>
<input>
<ID>IN_0</ID>287 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add5</lparam></gate>
<gate>
<ID>185</ID>
<type>DE_TO</type>
<position>105.5,-20</position>
<input>
<ID>IN_0</ID>73 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr5</lparam></gate>
<gate>
<ID>57</ID>
<type>DA_FROM</type>
<position>55,-32.5</position>
<input>
<ID>IN_0</ID>291 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr6</lparam></gate>
<gate>
<ID>187</ID>
<type>DE_TO</type>
<position>105.5,-22</position>
<input>
<ID>IN_0</ID>497 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr4</lparam></gate>
<gate>
<ID>59</ID>
<type>DE_TO</type>
<position>67,-38</position>
<input>
<ID>IN_0</ID>289 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add7</lparam></gate>
<gate>
<ID>747</ID>
<type>DE_TO</type>
<position>229,-115</position>
<input>
<ID>IN_0</ID>991 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN6</lparam></gate>
<gate>
<ID>61</ID>
<type>DA_FROM</type>
<position>55,-30.5</position>
<input>
<ID>IN_0</ID>290 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr5</lparam></gate>
<gate>
<ID>63</ID>
<type>DA_FROM</type>
<position>55,-37</position>
<input>
<ID>IN_0</ID>294 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac4</lparam></gate>
<gate>
<ID>64</ID>
<type>DA_FROM</type>
<position>55,-39</position>
<input>
<ID>IN_0</ID>295 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac5</lparam></gate>
<gate>
<ID>65</ID>
<type>DA_FROM</type>
<position>55,-41</position>
<input>
<ID>IN_0</ID>296 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac6</lparam></gate>
<gate>
<ID>67</ID>
<type>DA_FROM</type>
<position>55,-43</position>
<input>
<ID>IN_0</ID>297 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac7</lparam></gate>
<gate>
<ID>71</ID>
<type>AE_FULLADDER_4BIT</type>
<position>61,-52</position>
<input>
<ID>IN_0</ID>445 </input>
<input>
<ID>IN_1</ID>446 </input>
<input>
<ID>IN_2</ID>447 </input>
<input>
<ID>IN_3</ID>448 </input>
<input>
<ID>IN_B_0</ID>444 </input>
<input>
<ID>IN_B_1</ID>441 </input>
<input>
<ID>IN_B_2</ID>442 </input>
<input>
<ID>IN_B_3</ID>443 </input>
<output>
<ID>OUT_0</ID>298 </output>
<output>
<ID>OUT_1</ID>299 </output>
<output>
<ID>OUT_2</ID>439 </output>
<output>
<ID>OUT_3</ID>440 </output>
<input>
<ID>carry_in</ID>462 </input>
<output>
<ID>carry_out</ID>463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>72</ID>
<type>DA_FROM</type>
<position>55,-51.5</position>
<input>
<ID>IN_0</ID>443 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr11</lparam></gate>
<gate>
<ID>138</ID>
<type>AE_REGISTER8</type>
<position>98,-23.5</position>
<input>
<ID>IN_0</ID>478 </input>
<input>
<ID>IN_1</ID>479 </input>
<input>
<ID>IN_2</ID>480 </input>
<input>
<ID>IN_3</ID>481 </input>
<input>
<ID>IN_4</ID>485 </input>
<input>
<ID>IN_5</ID>484 </input>
<input>
<ID>IN_6</ID>483 </input>
<input>
<ID>IN_7</ID>482 </input>
<output>
<ID>OUT_0</ID>489 </output>
<output>
<ID>OUT_1</ID>496 </output>
<output>
<ID>OUT_2</ID>495 </output>
<output>
<ID>OUT_3</ID>494 </output>
<output>
<ID>OUT_4</ID>497 </output>
<output>
<ID>OUT_5</ID>73 </output>
<output>
<ID>OUT_6</ID>491 </output>
<output>
<ID>OUT_7</ID>490 </output>
<input>
<ID>clock</ID>488 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>74</ID>
<type>DA_FROM</type>
<position>55,-45.5</position>
<input>
<ID>IN_0</ID>444 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr8</lparam></gate>
<gate>
<ID>76</ID>
<type>DA_FROM</type>
<position>55,-49.5</position>
<input>
<ID>IN_0</ID>442 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr10</lparam></gate>
<gate>
<ID>78</ID>
<type>DA_FROM</type>
<position>55,-47.5</position>
<input>
<ID>IN_0</ID>441 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr9</lparam></gate>
<gate>
<ID>79</ID>
<type>DA_FROM</type>
<position>55,-54</position>
<input>
<ID>IN_0</ID>445 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac8</lparam></gate>
<gate>
<ID>81</ID>
<type>DA_FROM</type>
<position>55,-58</position>
<input>
<ID>IN_0</ID>447 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac10</lparam></gate>
<gate>
<ID>82</ID>
<type>DA_FROM</type>
<position>55,-60</position>
<input>
<ID>IN_0</ID>448 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac11</lparam></gate>
<gate>
<ID>83</ID>
<type>DE_TO</type>
<position>67,-70</position>
<input>
<ID>IN_0</ID>451 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add14</lparam></gate>
<gate>
<ID>85</ID>
<type>DA_FROM</type>
<position>55,-68.5</position>
<input>
<ID>IN_0</ID>455 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr15</lparam></gate>
<gate>
<ID>86</ID>
<type>DE_TO</type>
<position>67,-66</position>
<input>
<ID>IN_0</ID>449 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add12</lparam></gate>
<gate>
<ID>87</ID>
<type>DA_FROM</type>
<position>55,-62.5</position>
<input>
<ID>IN_0</ID>456 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr12</lparam></gate>
<gate>
<ID>168</ID>
<type>DE_TO</type>
<position>105.5,-18</position>
<input>
<ID>IN_0</ID>491 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr6</lparam></gate>
<gate>
<ID>471</ID>
<type>DA_FROM</type>
<position>140,-152.5</position>
<input>
<ID>IN_0</ID>710 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR</lparam></gate>
<gate>
<ID>104</ID>
<type>DE_TO</type>
<position>67,-68</position>
<input>
<ID>IN_0</ID>450 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add13</lparam></gate>
<gate>
<ID>465</ID>
<type>AA_AND2</type>
<position>145,-177.5</position>
<input>
<ID>IN_0</ID>719 </input>
<input>
<ID>IN_1</ID>938 </input>
<output>
<ID>OUT</ID>725 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>106</ID>
<type>DA_FROM</type>
<position>55,-66.5</position>
<input>
<ID>IN_0</ID>454 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr14</lparam></gate>
<gate>
<ID>108</ID>
<type>DE_TO</type>
<position>67,-72</position>
<input>
<ID>IN_0</ID>452 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add15</lparam></gate>
<gate>
<ID>459</ID>
<type>AA_AND2</type>
<position>197,-153.5</position>
<input>
<ID>IN_0</ID>734 </input>
<input>
<ID>IN_1</ID>942 </input>
<output>
<ID>OUT</ID>747 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>110</ID>
<type>DA_FROM</type>
<position>55,-64.5</position>
<input>
<ID>IN_0</ID>453 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr13</lparam></gate>
<gate>
<ID>469</ID>
<type>DA_FROM</type>
<position>140,-146.5</position>
<input>
<ID>IN_0</ID>708 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>479</ID>
<type>DE_TO</type>
<position>117.5,-26</position>
<input>
<ID>IN_0</ID>608 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr13</lparam></gate>
<gate>
<ID>112</ID>
<type>DA_FROM</type>
<position>55,-71</position>
<input>
<ID>IN_0</ID>457 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac12</lparam></gate>
<gate>
<ID>114</ID>
<type>DA_FROM</type>
<position>55,-73</position>
<input>
<ID>IN_0</ID>458 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac13</lparam></gate>
<gate>
<ID>473</ID>
<type>DA_FROM</type>
<position>140,-158.5</position>
<input>
<ID>IN_0</ID>712 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>116</ID>
<type>DA_FROM</type>
<position>55,-75</position>
<input>
<ID>IN_0</ID>459 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac14</lparam></gate>
<gate>
<ID>122</ID>
<type>DE_TO</type>
<position>60,-79</position>
<input>
<ID>IN_0</ID>464 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Cout</lparam></gate>
<gate>
<ID>481</ID>
<type>DE_OR8</type>
<position>170.5,-160</position>
<input>
<ID>IN_0</ID>721 </input>
<input>
<ID>IN_1</ID>722 </input>
<input>
<ID>IN_2</ID>723 </input>
<input>
<ID>IN_3</ID>724 </input>
<input>
<ID>IN_4</ID>331 </input>
<input>
<ID>IN_5</ID>725 </input>
<input>
<ID>IN_6</ID>726 </input>
<input>
<ID>IN_7</ID>727 </input>
<output>
<ID>OUT</ID>994 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>126</ID>
<type>FF_GND</type>
<position>66,-11</position>
<output>
<ID>OUT_0</ID>465 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>485</ID>
<type>AA_AND2</type>
<position>197,-159.5</position>
<input>
<ID>IN_0</ID>736 </input>
<input>
<ID>IN_1</ID>943 </input>
<output>
<ID>OUT</ID>748 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>130</ID>
<type>DD_KEYPAD_HEX</type>
<position>85.5,-17</position>
<output>
<ID>OUT_0</ID>485 </output>
<output>
<ID>OUT_1</ID>484 </output>
<output>
<ID>OUT_2</ID>483 </output>
<output>
<ID>OUT_3</ID>482 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>134</ID>
<type>DD_KEYPAD_HEX</type>
<position>85.5,-29</position>
<output>
<ID>OUT_0</ID>478 </output>
<output>
<ID>OUT_1</ID>479 </output>
<output>
<ID>OUT_2</ID>480 </output>
<output>
<ID>OUT_3</ID>481 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>158</ID>
<type>DA_FROM</type>
<position>97,-30.5</position>
<input>
<ID>IN_0</ID>488 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>162</ID>
<type>DE_TO</type>
<position>105.5,-30</position>
<input>
<ID>IN_0</ID>489 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr0</lparam></gate>
<gate>
<ID>166</ID>
<type>DE_TO</type>
<position>105.5,-16</position>
<input>
<ID>IN_0</ID>490 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr7</lparam></gate>
<gate>
<ID>219</ID>
<type>DE_TO</type>
<position>105.5,-24</position>
<input>
<ID>IN_0</ID>494 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr3</lparam></gate>
<gate>
<ID>380</ID>
<type>AA_AND2</type>
<position>197.5,-114.5</position>
<input>
<ID>IN_0</ID>640 </input>
<input>
<ID>IN_1</ID>911 </input>
<output>
<ID>OUT</ID>652 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>557</ID>
<type>AA_AND3</type>
<position>145,-186</position>
<input>
<ID>IN_0</ID>801 </input>
<input>
<ID>IN_1</ID>963 </input>
<input>
<ID>IN_2</ID>964 </input>
<output>
<ID>OUT</ID>817 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>220</ID>
<type>DE_TO</type>
<position>105.5,-26</position>
<input>
<ID>IN_0</ID>495 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr2</lparam></gate>
<gate>
<ID>550</ID>
<type>DA_FROM</type>
<position>88.5,-216</position>
<input>
<ID>IN_0</ID>789 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>221</ID>
<type>DE_TO</type>
<position>105.5,-28</position>
<input>
<ID>IN_0</ID>496 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr1</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_AND3</type>
<position>94,-50</position>
<input>
<ID>IN_0</ID>466 </input>
<input>
<ID>IN_1</ID>467 </input>
<input>
<ID>IN_2</ID>468 </input>
<output>
<ID>OUT</ID>501 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_AND2</type>
<position>94,-57</position>
<input>
<ID>IN_0</ID>469 </input>
<input>
<ID>IN_1</ID>470 </input>
<output>
<ID>OUT</ID>502 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>120</ID>
<type>AA_AND2</type>
<position>94,-63</position>
<input>
<ID>IN_0</ID>473 </input>
<input>
<ID>IN_1</ID>474 </input>
<output>
<ID>OUT</ID>503 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>487</ID>
<type>AA_AND2</type>
<position>197,-171.5</position>
<input>
<ID>IN_0</ID>741 </input>
<input>
<ID>IN_1</ID>945 </input>
<output>
<ID>OUT</ID>750 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>124</ID>
<type>AA_AND2</type>
<position>94,-69</position>
<input>
<ID>IN_0</ID>475 </input>
<input>
<ID>IN_1</ID>476 </input>
<output>
<ID>OUT</ID>508 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>475</ID>
<type>DA_FROM</type>
<position>140,-164.5</position>
<input>
<ID>IN_0</ID>714 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>128</ID>
<type>AA_AND2</type>
<position>94,-75</position>
<input>
<ID>IN_0</ID>477 </input>
<input>
<ID>IN_1</ID>487 </input>
<output>
<ID>OUT</ID>511 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>132</ID>
<type>AA_AND2</type>
<position>94,-81</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>498 </input>
<output>
<ID>OUT</ID>510 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>136</ID>
<type>AA_AND2</type>
<position>94,-87</position>
<input>
<ID>IN_0</ID>499 </input>
<input>
<ID>IN_1</ID>348 </input>
<output>
<ID>OUT</ID>509 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>142</ID>
<type>DA_FROM</type>
<position>89,-48</position>
<input>
<ID>IN_0</ID>466 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>146</ID>
<type>DA_FROM</type>
<position>89,-50</position>
<input>
<ID>IN_0</ID>467 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr0</lparam></gate>
<gate>
<ID>150</ID>
<type>DA_FROM</type>
<position>89,-52</position>
<input>
<ID>IN_0</ID>468 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac0</lparam></gate>
<gate>
<ID>154</ID>
<type>DA_FROM</type>
<position>89,-56</position>
<input>
<ID>IN_0</ID>469 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>160</ID>
<type>DA_FROM</type>
<position>89,-58</position>
<input>
<ID>IN_0</ID>470 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add0</lparam></gate>
<gate>
<ID>226</ID>
<type>DA_FROM</type>
<position>89,-62</position>
<input>
<ID>IN_0</ID>473 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR</lparam></gate>
<gate>
<ID>228</ID>
<type>DA_FROM</type>
<position>89,-64</position>
<input>
<ID>IN_0</ID>474 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr0</lparam></gate>
<gate>
<ID>558</ID>
<type>AA_AND2</type>
<position>145,-193</position>
<input>
<ID>IN_0</ID>804 </input>
<input>
<ID>IN_1</ID>965 </input>
<output>
<ID>OUT</ID>818 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>230</ID>
<type>DA_FROM</type>
<position>89,-68</position>
<input>
<ID>IN_0</ID>475 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>232</ID>
<type>DA_FROM</type>
<position>89,-70</position>
<input>
<ID>IN_0</ID>476 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr0</lparam></gate>
<gate>
<ID>562</ID>
<type>DA_FROM</type>
<position>140,-222</position>
<input>
<ID>IN_0</ID>815 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>234</ID>
<type>DA_FROM</type>
<position>89,-74</position>
<input>
<ID>IN_0</ID>477 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>236</ID>
<type>DA_FROM</type>
<position>85,-76</position>
<input>
<ID>IN_0</ID>492 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac0</lparam></gate>
<gate>
<ID>566</ID>
<type>DA_FROM</type>
<position>140,-184</position>
<input>
<ID>IN_0</ID>801 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>238</ID>
<type>AE_SMALL_INVERTER</type>
<position>89,-76</position>
<input>
<ID>IN_0</ID>492 </input>
<output>
<ID>OUT_0</ID>487 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>240</ID>
<type>DA_FROM</type>
<position>89,-80</position>
<input>
<ID>IN_0</ID>493 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>242</ID>
<type>DA_FROM</type>
<position>89,-82</position>
<input>
<ID>IN_0</ID>498 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac1</lparam></gate>
<gate>
<ID>244</ID>
<type>DA_FROM</type>
<position>89,-86</position>
<input>
<ID>IN_0</ID>499 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>248</ID>
<type>DE_OR8</type>
<position>119.5,-69.5</position>
<input>
<ID>IN_0</ID>501 </input>
<input>
<ID>IN_1</ID>502 </input>
<input>
<ID>IN_2</ID>503 </input>
<input>
<ID>IN_3</ID>508 </input>
<input>
<ID>IN_4</ID>536 </input>
<input>
<ID>IN_5</ID>509 </input>
<input>
<ID>IN_6</ID>510 </input>
<input>
<ID>IN_7</ID>511 </input>
<output>
<ID>OUT</ID>512 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>250</ID>
<type>DE_TO</type>
<position>125.5,-69.5</position>
<input>
<ID>IN_0</ID>512 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN0</lparam></gate>
<gate>
<ID>251</ID>
<type>AA_AND3</type>
<position>145.5,-50</position>
<input>
<ID>IN_0</ID>513 </input>
<input>
<ID>IN_1</ID>514 </input>
<input>
<ID>IN_2</ID>515 </input>
<output>
<ID>OUT</ID>529 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>252</ID>
<type>AA_AND2</type>
<position>145.5,-57</position>
<input>
<ID>IN_0</ID>516 </input>
<input>
<ID>IN_1</ID>517 </input>
<output>
<ID>OUT</ID>530 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>253</ID>
<type>AA_AND2</type>
<position>145.5,-63</position>
<input>
<ID>IN_0</ID>518 </input>
<input>
<ID>IN_1</ID>519 </input>
<output>
<ID>OUT</ID>531 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>278</ID>
<type>AA_AND2</type>
<position>197.5,-63</position>
<input>
<ID>IN_0</ID>542 </input>
<input>
<ID>IN_1</ID>877 </input>
<output>
<ID>OUT</ID>555 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>254</ID>
<type>AA_AND2</type>
<position>145.5,-69</position>
<input>
<ID>IN_0</ID>520 </input>
<input>
<ID>IN_1</ID>521 </input>
<output>
<ID>OUT</ID>532 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>255</ID>
<type>AA_AND2</type>
<position>145.5,-75</position>
<input>
<ID>IN_0</ID>522 </input>
<input>
<ID>IN_1</ID>523 </input>
<output>
<ID>OUT</ID>535 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>272</ID>
<type>DA_FROM</type>
<position>140.5,-86</position>
<input>
<ID>IN_0</ID>527 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>256</ID>
<type>AA_AND2</type>
<position>145.5,-81</position>
<input>
<ID>IN_0</ID>525 </input>
<input>
<ID>IN_1</ID>526 </input>
<output>
<ID>OUT</ID>534 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>561</ID>
<type>AA_AND2</type>
<position>145,-205</position>
<input>
<ID>IN_0</ID>808 </input>
<input>
<ID>IN_1</ID>967 </input>
<output>
<ID>OUT</ID>820 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>239</ID>
<type>FF_GND</type>
<position>116.5,-74.5</position>
<output>
<ID>OUT_0</ID>536 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>257</ID>
<type>AA_AND2</type>
<position>145.5,-87</position>
<input>
<ID>IN_0</ID>527 </input>
<input>
<ID>IN_1</ID>881 </input>
<output>
<ID>OUT</ID>533 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>592</ID>
<type>DA_FROM</type>
<position>192,-204</position>
<input>
<ID>IN_0</ID>832 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>258</ID>
<type>DA_FROM</type>
<position>140.5,-48</position>
<input>
<ID>IN_0</ID>513 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>233</ID>
<type>FF_GND</type>
<position>271.5,-74.5</position>
<output>
<ID>OUT_0</ID>506 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>259</ID>
<type>DA_FROM</type>
<position>140.5,-50</position>
<input>
<ID>IN_0</ID>514 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr1</lparam></gate>
<gate>
<ID>750</ID>
<type>DE_TO</type>
<position>176.5,-160</position>
<input>
<ID>IN_0</ID>994 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN9</lparam></gate>
<gate>
<ID>260</ID>
<type>DA_FROM</type>
<position>140.5,-52</position>
<input>
<ID>IN_0</ID>515 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac1</lparam></gate>
<gate>
<ID>565</ID>
<type>AA_AND2</type>
<position>145,-223</position>
<input>
<ID>IN_0</ID>815 </input>
<input>
<ID>IN_1</ID>970 </input>
<output>
<ID>OUT</ID>821 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>227</ID>
<type>FF_GND</type>
<position>220,-120</position>
<output>
<ID>OUT_0</ID>500 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>261</ID>
<type>DA_FROM</type>
<position>140.5,-56</position>
<input>
<ID>IN_0</ID>516 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>596</ID>
<type>DA_FROM</type>
<position>192,-216</position>
<input>
<ID>IN_0</ID>837 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>262</ID>
<type>DA_FROM</type>
<position>140.5,-58</position>
<input>
<ID>IN_0</ID>517 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add1</lparam></gate>
<gate>
<ID>237</ID>
<type>FF_GND</type>
<position>168,-74.5</position>
<output>
<ID>OUT_0</ID>528 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>263</ID>
<type>DA_FROM</type>
<position>140.5,-62</position>
<input>
<ID>IN_0</ID>518 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR</lparam></gate>
<gate>
<ID>738</ID>
<type>DA_FROM</type>
<position>243.5,-200</position>
<input>
<ID>IN_0</ID>982 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr15</lparam></gate>
<gate>
<ID>264</ID>
<type>DA_FROM</type>
<position>140.5,-64</position>
<input>
<ID>IN_0</ID>519 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr1</lparam></gate>
<gate>
<ID>569</ID>
<type>DA_FROM</type>
<position>140,-192</position>
<input>
<ID>IN_0</ID>804 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>265</ID>
<type>DA_FROM</type>
<position>140.5,-68</position>
<input>
<ID>IN_0</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>600</ID>
<type>DE_OR8</type>
<position>222.5,-205.5</position>
<input>
<ID>IN_0</ID>841 </input>
<input>
<ID>IN_1</ID>842 </input>
<input>
<ID>IN_2</ID>843 </input>
<input>
<ID>IN_3</ID>844 </input>
<input>
<ID>IN_4</ID>104 </input>
<input>
<ID>IN_5</ID>845 </input>
<input>
<ID>IN_6</ID>846 </input>
<input>
<ID>IN_7</ID>847 </input>
<output>
<ID>OUT</ID>999 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>266</ID>
<type>DA_FROM</type>
<position>140.5,-70</position>
<input>
<ID>IN_0</ID>521 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr1</lparam></gate>
<gate>
<ID>267</ID>
<type>DA_FROM</type>
<position>140.5,-74</position>
<input>
<ID>IN_0</ID>522 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>268</ID>
<type>DA_FROM</type>
<position>136.5,-76</position>
<input>
<ID>IN_0</ID>524 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac1</lparam></gate>
<gate>
<ID>573</ID>
<type>DA_FROM</type>
<position>140,-204</position>
<input>
<ID>IN_0</ID>808 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>235</ID>
<type>FF_GND</type>
<position>220,-74.5</position>
<output>
<ID>OUT_0</ID>507 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>269</ID>
<type>AE_SMALL_INVERTER</type>
<position>140.5,-76</position>
<input>
<ID>IN_0</ID>524 </input>
<output>
<ID>OUT_0</ID>523 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>604</ID>
<type>AA_AND2</type>
<position>248.5,-199</position>
<input>
<ID>IN_0</ID>854 </input>
<input>
<ID>IN_1</ID>982 </input>
<output>
<ID>OUT</ID>867 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>270</ID>
<type>DA_FROM</type>
<position>140.5,-80</position>
<input>
<ID>IN_0</ID>525 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>271</ID>
<type>DA_FROM</type>
<position>140.5,-82</position>
<input>
<ID>IN_0</ID>526 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac2</lparam></gate>
<gate>
<ID>746</ID>
<type>DE_TO</type>
<position>177,-115</position>
<input>
<ID>IN_0</ID>990 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN5</lparam></gate>
<gate>
<ID>608</ID>
<type>AA_AND2</type>
<position>248.5,-217</position>
<input>
<ID>IN_0</ID>861 </input>
<input>
<ID>IN_1</ID>862 </input>
<output>
<ID>OUT</ID>870 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>274</ID>
<type>DE_OR8</type>
<position>171,-69.5</position>
<input>
<ID>IN_0</ID>529 </input>
<input>
<ID>IN_1</ID>530 </input>
<input>
<ID>IN_2</ID>531 </input>
<input>
<ID>IN_3</ID>532 </input>
<input>
<ID>IN_4</ID>528 </input>
<input>
<ID>IN_5</ID>533 </input>
<input>
<ID>IN_6</ID>534 </input>
<input>
<ID>IN_7</ID>535 </input>
<output>
<ID>OUT</ID>986 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>276</ID>
<type>AA_AND3</type>
<position>197.5,-50</position>
<input>
<ID>IN_0</ID>537 </input>
<input>
<ID>IN_1</ID>874 </input>
<input>
<ID>IN_2</ID>875 </input>
<output>
<ID>OUT</ID>553 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>243</ID>
<type>FF_GND</type>
<position>90,-89</position>
<output>
<ID>OUT_0</ID>348 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>277</ID>
<type>AA_AND2</type>
<position>197.5,-57</position>
<input>
<ID>IN_0</ID>540 </input>
<input>
<ID>IN_1</ID>876 </input>
<output>
<ID>OUT</ID>554 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>279</ID>
<type>AA_AND2</type>
<position>197.5,-69</position>
<input>
<ID>IN_0</ID>544 </input>
<input>
<ID>IN_1</ID>878 </input>
<output>
<ID>OUT</ID>556 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>754</ID>
<type>DE_TO</type>
<position>176.5,-205.5</position>
<input>
<ID>IN_0</ID>998 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN13</lparam></gate>
<gate>
<ID>280</ID>
<type>AA_AND2</type>
<position>197.5,-75</position>
<input>
<ID>IN_0</ID>546 </input>
<input>
<ID>IN_1</ID>547 </input>
<output>
<ID>OUT</ID>559 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>281</ID>
<type>AA_AND2</type>
<position>197.5,-81</position>
<input>
<ID>IN_0</ID>549 </input>
<input>
<ID>IN_1</ID>880 </input>
<output>
<ID>OUT</ID>558 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>616</ID>
<type>DA_FROM</type>
<position>243.5,-204</position>
<input>
<ID>IN_0</ID>856 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>282</ID>
<type>AA_AND2</type>
<position>197.5,-87</position>
<input>
<ID>IN_0</ID>551 </input>
<input>
<ID>IN_1</ID>882 </input>
<output>
<ID>OUT</ID>557 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>283</ID>
<type>DA_FROM</type>
<position>192.5,-48</position>
<input>
<ID>IN_0</ID>537 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>646</ID>
<type>DA_FROM</type>
<position>89,-103.5</position>
<input>
<ID>IN_0</ID>893 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add4</lparam></gate>
<gate>
<ID>620</ID>
<type>AE_SMALL_INVERTER</type>
<position>243.5,-212</position>
<input>
<ID>IN_0</ID>984 </input>
<output>
<ID>OUT_0</ID>859 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>286</ID>
<type>DA_FROM</type>
<position>192.5,-56</position>
<input>
<ID>IN_0</ID>540 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>288</ID>
<type>DA_FROM</type>
<position>192.5,-62</position>
<input>
<ID>IN_0</ID>542 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR</lparam></gate>
<gate>
<ID>624</ID>
<type>DE_OR8</type>
<position>274,-205.5</position>
<input>
<ID>IN_0</ID>865 </input>
<input>
<ID>IN_1</ID>866 </input>
<input>
<ID>IN_2</ID>867 </input>
<input>
<ID>IN_3</ID>868 </input>
<input>
<ID>IN_4</ID>97 </input>
<input>
<ID>IN_5</ID>869 </input>
<input>
<ID>IN_6</ID>870 </input>
<input>
<ID>IN_7</ID>871 </input>
<output>
<ID>OUT</ID>1000 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>290</ID>
<type>DA_FROM</type>
<position>192.5,-68</position>
<input>
<ID>IN_0</ID>544 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>292</ID>
<type>DA_FROM</type>
<position>192.5,-74</position>
<input>
<ID>IN_0</ID>546 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>628</ID>
<type>DA_FROM</type>
<position>192.5,-52</position>
<input>
<ID>IN_0</ID>875 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac2</lparam></gate>
<gate>
<ID>294</ID>
<type>AE_SMALL_INVERTER</type>
<position>192.5,-76</position>
<input>
<ID>IN_0</ID>879 </input>
<output>
<ID>OUT_0</ID>547 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>295</ID>
<type>DA_FROM</type>
<position>192.5,-80</position>
<input>
<ID>IN_0</ID>549 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>642</ID>
<type>DA_FROM</type>
<position>244,-82</position>
<input>
<ID>IN_0</ID>889 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac4</lparam></gate>
<gate>
<ID>297</ID>
<type>DA_FROM</type>
<position>192.5,-86</position>
<input>
<ID>IN_0</ID>551 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>632</ID>
<type>DA_FROM</type>
<position>188.5,-76</position>
<input>
<ID>IN_0</ID>879 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac2</lparam></gate>
<gate>
<ID>299</ID>
<type>DE_OR8</type>
<position>223,-69.5</position>
<input>
<ID>IN_0</ID>553 </input>
<input>
<ID>IN_1</ID>554 </input>
<input>
<ID>IN_2</ID>555 </input>
<input>
<ID>IN_3</ID>556 </input>
<input>
<ID>IN_4</ID>507 </input>
<input>
<ID>IN_5</ID>557 </input>
<input>
<ID>IN_6</ID>558 </input>
<input>
<ID>IN_7</ID>559 </input>
<output>
<ID>OUT</ID>987 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>662</ID>
<type>DA_FROM</type>
<position>192.5,-103.5</position>
<input>
<ID>IN_0</ID>909 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add6</lparam></gate>
<gate>
<ID>301</ID>
<type>AA_AND3</type>
<position>249,-50</position>
<input>
<ID>IN_0</ID>561 </input>
<input>
<ID>IN_1</ID>883 </input>
<input>
<ID>IN_2</ID>884 </input>
<output>
<ID>OUT</ID>577 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>636</ID>
<type>DA_FROM</type>
<position>244,-50</position>
<input>
<ID>IN_0</ID>883 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr3</lparam></gate>
<gate>
<ID>302</ID>
<type>AA_AND2</type>
<position>249,-57</position>
<input>
<ID>IN_0</ID>564 </input>
<input>
<ID>IN_1</ID>885 </input>
<output>
<ID>OUT</ID>578 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>303</ID>
<type>AA_AND2</type>
<position>249,-63</position>
<input>
<ID>IN_0</ID>566 </input>
<input>
<ID>IN_1</ID>886 </input>
<output>
<ID>OUT</ID>579 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>650</ID>
<type>DA_FROM</type>
<position>89,-127.5</position>
<input>
<ID>IN_0</ID>897 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac5</lparam></gate>
<gate>
<ID>304</ID>
<type>AA_AND2</type>
<position>249,-69</position>
<input>
<ID>IN_0</ID>568 </input>
<input>
<ID>IN_1</ID>887 </input>
<output>
<ID>OUT</ID>580 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>305</ID>
<type>DA_FROM</type>
<position>244,-86</position>
<input>
<ID>IN_0</ID>575 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>512</ID>
<type>AA_AND2</type>
<position>248.5,-171.5</position>
<input>
<ID>IN_0</ID>765 </input>
<input>
<ID>IN_1</ID>953 </input>
<output>
<ID>OUT</ID>774 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>306</ID>
<type>AA_AND2</type>
<position>249,-75</position>
<input>
<ID>IN_0</ID>570 </input>
<input>
<ID>IN_1</ID>571 </input>
<output>
<ID>OUT</ID>583 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>307</ID>
<type>AA_AND2</type>
<position>249,-81</position>
<input>
<ID>IN_0</ID>573 </input>
<input>
<ID>IN_1</ID>889 </input>
<output>
<ID>OUT</ID>582 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>670</ID>
<type>DA_FROM</type>
<position>244,-103.5</position>
<input>
<ID>IN_0</ID>917 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add7</lparam></gate>
<gate>
<ID>308</ID>
<type>AA_AND2</type>
<position>249,-87</position>
<input>
<ID>IN_0</ID>575 </input>
<input>
<ID>IN_1</ID>890 </input>
<output>
<ID>OUT</ID>581 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>309</ID>
<type>DA_FROM</type>
<position>244,-48</position>
<input>
<ID>IN_0</ID>561 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>312</ID>
<type>DA_FROM</type>
<position>244,-56</position>
<input>
<ID>IN_0</ID>564 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>314</ID>
<type>DA_FROM</type>
<position>244,-62</position>
<input>
<ID>IN_0</ID>566 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR</lparam></gate>
<gate>
<ID>316</ID>
<type>DA_FROM</type>
<position>244,-68</position>
<input>
<ID>IN_0</ID>568 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>318</ID>
<type>DA_FROM</type>
<position>244,-74</position>
<input>
<ID>IN_0</ID>570 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>320</ID>
<type>AE_SMALL_INVERTER</type>
<position>244,-76</position>
<input>
<ID>IN_0</ID>888 </input>
<output>
<ID>OUT_0</ID>571 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>321</ID>
<type>DA_FROM</type>
<position>244,-80</position>
<input>
<ID>IN_0</ID>573 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>656</ID>
<type>DA_FROM</type>
<position>140.5,-115.5</position>
<input>
<ID>IN_0</ID>903 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr5</lparam></gate>
<gate>
<ID>324</ID>
<type>DE_OR8</type>
<position>274.5,-69.5</position>
<input>
<ID>IN_0</ID>577 </input>
<input>
<ID>IN_1</ID>578 </input>
<input>
<ID>IN_2</ID>579 </input>
<input>
<ID>IN_3</ID>580 </input>
<input>
<ID>IN_4</ID>506 </input>
<input>
<ID>IN_5</ID>581 </input>
<input>
<ID>IN_6</ID>582 </input>
<input>
<ID>IN_7</ID>583 </input>
<output>
<ID>OUT</ID>988 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>629</ID>
<type>DA_FROM</type>
<position>192.5,-58</position>
<input>
<ID>IN_0</ID>876 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add2</lparam></gate>
<gate>
<ID>660</ID>
<type>DA_FROM</type>
<position>192.5,-95.5</position>
<input>
<ID>IN_0</ID>907 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr6</lparam></gate>
<gate>
<ID>326</ID>
<type>AA_AND3</type>
<position>94,-95.5</position>
<input>
<ID>IN_0</ID>585 </input>
<input>
<ID>IN_1</ID>891 </input>
<input>
<ID>IN_2</ID>892 </input>
<output>
<ID>OUT</ID>601 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>327</ID>
<type>AA_AND2</type>
<position>94,-102.5</position>
<input>
<ID>IN_0</ID>588 </input>
<input>
<ID>IN_1</ID>893 </input>
<output>
<ID>OUT</ID>602 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>328</ID>
<type>AA_AND2</type>
<position>94,-108.5</position>
<input>
<ID>IN_0</ID>590 </input>
<input>
<ID>IN_1</ID>894 </input>
<output>
<ID>OUT</ID>603 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>633</ID>
<type>DA_FROM</type>
<position>192.5,-82</position>
<input>
<ID>IN_0</ID>880 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac3</lparam></gate>
<gate>
<ID>329</ID>
<type>AA_AND2</type>
<position>94,-114.5</position>
<input>
<ID>IN_0</ID>592 </input>
<input>
<ID>IN_1</ID>895 </input>
<output>
<ID>OUT</ID>604 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>664</ID>
<type>DA_FROM</type>
<position>192.5,-115.5</position>
<input>
<ID>IN_0</ID>911 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr6</lparam></gate>
<gate>
<ID>330</ID>
<type>AA_AND2</type>
<position>94,-120.5</position>
<input>
<ID>IN_0</ID>594 </input>
<input>
<ID>IN_1</ID>595 </input>
<output>
<ID>OUT</ID>607 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>331</ID>
<type>AA_AND2</type>
<position>94,-126.5</position>
<input>
<ID>IN_0</ID>597 </input>
<input>
<ID>IN_1</ID>897 </input>
<output>
<ID>OUT</ID>606 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>332</ID>
<type>AA_AND2</type>
<position>94,-132.5</position>
<input>
<ID>IN_0</ID>599 </input>
<input>
<ID>IN_1</ID>898 </input>
<output>
<ID>OUT</ID>605 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>637</ID>
<type>DA_FROM</type>
<position>244,-52</position>
<input>
<ID>IN_0</ID>884 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac3</lparam></gate>
<gate>
<ID>333</ID>
<type>DA_FROM</type>
<position>89,-93.5</position>
<input>
<ID>IN_0</ID>585 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>668</ID>
<type>DA_FROM</type>
<position>244,-95.5</position>
<input>
<ID>IN_0</ID>915 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr7</lparam></gate>
<gate>
<ID>336</ID>
<type>DA_FROM</type>
<position>89,-101.5</position>
<input>
<ID>IN_0</ID>588 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>513</ID>
<type>AA_AND2</type>
<position>248.5,-177.5</position>
<input>
<ID>IN_0</ID>767 </input>
<input>
<ID>IN_1</ID>954 </input>
<output>
<ID>OUT</ID>773 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>338</ID>
<type>DA_FROM</type>
<position>89,-107.5</position>
<input>
<ID>IN_0</ID>590 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR</lparam></gate>
<gate>
<ID>340</ID>
<type>DA_FROM</type>
<position>89,-113.5</position>
<input>
<ID>IN_0</ID>592 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>517</ID>
<type>DA_FROM</type>
<position>243.5,-146.5</position>
<input>
<ID>IN_0</ID>756 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>342</ID>
<type>DA_FROM</type>
<position>89,-119.5</position>
<input>
<ID>IN_0</ID>594 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>344</ID>
<type>AE_SMALL_INVERTER</type>
<position>89,-121.5</position>
<input>
<ID>IN_0</ID>896 </input>
<output>
<ID>OUT_0</ID>595 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>521</ID>
<type>DA_FROM</type>
<position>243.5,-158.5</position>
<input>
<ID>IN_0</ID>760 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>345</ID>
<type>DA_FROM</type>
<position>89,-125.5</position>
<input>
<ID>IN_0</ID>597 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>680</ID>
<type>DA_FROM</type>
<position>88.5,-160.5</position>
<input>
<ID>IN_0</ID>927 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr8</lparam></gate>
<gate>
<ID>347</ID>
<type>DA_FROM</type>
<position>89,-131.5</position>
<input>
<ID>IN_0</ID>599 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>710</ID>
<type>DA_FROM</type>
<position>243.5,-178.5</position>
<input>
<ID>IN_0</ID>954 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac10</lparam></gate>
<gate>
<ID>525</ID>
<type>AE_SMALL_INVERTER</type>
<position>243.5,-166.5</position>
<input>
<ID>IN_0</ID>952 </input>
<output>
<ID>OUT_0</ID>763 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>349</ID>
<type>DE_OR8</type>
<position>119.5,-115</position>
<input>
<ID>IN_0</ID>601 </input>
<input>
<ID>IN_1</ID>602 </input>
<input>
<ID>IN_2</ID>603 </input>
<input>
<ID>IN_3</ID>604 </input>
<input>
<ID>IN_4</ID>505 </input>
<input>
<ID>IN_5</ID>605 </input>
<input>
<ID>IN_6</ID>606 </input>
<input>
<ID>IN_7</ID>607 </input>
<output>
<ID>OUT</ID>989 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>352</ID>
<type>AA_AND3</type>
<position>145.5,-95.5</position>
<input>
<ID>IN_0</ID>609 </input>
<input>
<ID>IN_1</ID>899 </input>
<input>
<ID>IN_2</ID>900 </input>
<output>
<ID>OUT</ID>625 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>529</ID>
<type>DE_OR8</type>
<position>274,-160</position>
<input>
<ID>IN_0</ID>769 </input>
<input>
<ID>IN_1</ID>770 </input>
<input>
<ID>IN_2</ID>771 </input>
<input>
<ID>IN_3</ID>772 </input>
<input>
<ID>IN_4</ID>472 </input>
<input>
<ID>IN_5</ID>773 </input>
<input>
<ID>IN_6</ID>774 </input>
<input>
<ID>IN_7</ID>775 </input>
<output>
<ID>OUT</ID>996 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>353</ID>
<type>AA_AND2</type>
<position>145.5,-102.5</position>
<input>
<ID>IN_0</ID>612 </input>
<input>
<ID>IN_1</ID>901 </input>
<output>
<ID>OUT</ID>626 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>688</ID>
<type>DA_FROM</type>
<position>140,-148.5</position>
<input>
<ID>IN_0</ID>933 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add9</lparam></gate>
<gate>
<ID>354</ID>
<type>AA_AND2</type>
<position>197.5,-108.5</position>
<input>
<ID>IN_0</ID>638 </input>
<input>
<ID>IN_1</ID>910 </input>
<output>
<ID>OUT</ID>651 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>355</ID>
<type>AA_AND2</type>
<position>145.5,-108.5</position>
<input>
<ID>IN_0</ID>614 </input>
<input>
<ID>IN_1</ID>902 </input>
<output>
<ID>OUT</ID>627 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>718</ID>
<type>DA_FROM</type>
<position>88.5,-224</position>
<input>
<ID>IN_0</ID>962 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac11</lparam></gate>
<gate>
<ID>356</ID>
<type>AA_AND2</type>
<position>145.5,-114.5</position>
<input>
<ID>IN_0</ID>616 </input>
<input>
<ID>IN_1</ID>903 </input>
<output>
<ID>OUT</ID>628 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>533</ID>
<type>AA_AND2</type>
<position>93.5,-199</position>
<input>
<ID>IN_0</ID>782 </input>
<input>
<ID>IN_1</ID>958 </input>
<output>
<ID>OUT</ID>795 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>357</ID>
<type>DA_FROM</type>
<position>140.5,-131.5</position>
<input>
<ID>IN_0</ID>623 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>692</ID>
<type>DA_FROM</type>
<position>140,-172.5</position>
<input>
<ID>IN_0</ID>937 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac10</lparam></gate>
<gate>
<ID>358</ID>
<type>AA_AND2</type>
<position>145.5,-120.5</position>
<input>
<ID>IN_0</ID>618 </input>
<input>
<ID>IN_1</ID>619 </input>
<output>
<ID>OUT</ID>631 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>359</ID>
<type>AA_AND2</type>
<position>145.5,-126.5</position>
<input>
<ID>IN_0</ID>621 </input>
<input>
<ID>IN_1</ID>905 </input>
<output>
<ID>OUT</ID>630 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>706</ID>
<type>DA_FROM</type>
<position>243.5,-154.5</position>
<input>
<ID>IN_0</ID>950 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr11</lparam></gate>
<gate>
<ID>360</ID>
<type>AA_AND2</type>
<position>145.5,-132.5</position>
<input>
<ID>IN_0</ID>623 </input>
<input>
<ID>IN_1</ID>906 </input>
<output>
<ID>OUT</ID>629 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>537</ID>
<type>AA_AND2</type>
<position>93.5,-223</position>
<input>
<ID>IN_0</ID>791 </input>
<input>
<ID>IN_1</ID>962 </input>
<output>
<ID>OUT</ID>797 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>361</ID>
<type>DA_FROM</type>
<position>140.5,-93.5</position>
<input>
<ID>IN_0</ID>609 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>696</ID>
<type>DA_FROM</type>
<position>192,-148.5</position>
<input>
<ID>IN_0</ID>941 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add10</lparam></gate>
<gate>
<ID>364</ID>
<type>DA_FROM</type>
<position>140.5,-101.5</position>
<input>
<ID>IN_0</ID>612 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>541</ID>
<type>DA_FROM</type>
<position>88.5,-192</position>
<input>
<ID>IN_0</ID>780 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>366</ID>
<type>DA_FROM</type>
<position>140.5,-107.5</position>
<input>
<ID>IN_0</ID>614 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR</lparam></gate>
<gate>
<ID>368</ID>
<type>DA_FROM</type>
<position>140.5,-113.5</position>
<input>
<ID>IN_0</ID>616 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>545</ID>
<type>DA_FROM</type>
<position>88.5,-204</position>
<input>
<ID>IN_0</ID>784 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>223</ID>
<type>FF_GND</type>
<position>219.5,-165</position>
<output>
<ID>OUT_0</ID>471 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>370</ID>
<type>DA_FROM</type>
<position>140.5,-119.5</position>
<input>
<ID>IN_0</ID>618 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>372</ID>
<type>AE_SMALL_INVERTER</type>
<position>140.5,-121.5</position>
<input>
<ID>IN_0</ID>904 </input>
<output>
<ID>OUT_0</ID>619 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>549</ID>
<type>AE_SMALL_INVERTER</type>
<position>88.5,-212</position>
<input>
<ID>IN_0</ID>960 </input>
<output>
<ID>OUT_0</ID>787 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>373</ID>
<type>DA_FROM</type>
<position>140.5,-125.5</position>
<input>
<ID>IN_0</ID>621 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>580</ID>
<type>DE_OR8</type>
<position>170.5,-205.5</position>
<input>
<ID>IN_0</ID>817 </input>
<input>
<ID>IN_1</ID>818 </input>
<input>
<ID>IN_2</ID>819 </input>
<input>
<ID>IN_3</ID>820 </input>
<input>
<ID>IN_4</ID>322 </input>
<input>
<ID>IN_5</ID>821 </input>
<input>
<ID>IN_6</ID>822 </input>
<input>
<ID>IN_7</ID>823 </input>
<output>
<ID>OUT</ID>998 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>376</ID>
<type>DE_OR8</type>
<position>171,-115</position>
<input>
<ID>IN_0</ID>625 </input>
<input>
<ID>IN_1</ID>626 </input>
<input>
<ID>IN_2</ID>627 </input>
<input>
<ID>IN_3</ID>628 </input>
<input>
<ID>IN_4</ID>504 </input>
<input>
<ID>IN_5</ID>629 </input>
<input>
<ID>IN_6</ID>630 </input>
<input>
<ID>IN_7</ID>631 </input>
<output>
<ID>OUT</ID>990 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>231</ID>
<type>FF_GND</type>
<position>116.5,-120</position>
<output>
<ID>OUT_0</ID>505 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>584</ID>
<type>AA_AND2</type>
<position>197,-211</position>
<input>
<ID>IN_0</ID>834 </input>
<input>
<ID>IN_1</ID>835 </input>
<output>
<ID>OUT</ID>847 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>378</ID>
<type>AA_AND3</type>
<position>197.5,-95.5</position>
<input>
<ID>IN_0</ID>633 </input>
<input>
<ID>IN_1</ID>907 </input>
<input>
<ID>IN_2</ID>908 </input>
<output>
<ID>OUT</ID>649 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>225</ID>
<type>FF_GND</type>
<position>271.5,-120</position>
<output>
<ID>OUT_0</ID>486 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>379</ID>
<type>AA_AND2</type>
<position>197.5,-102.5</position>
<input>
<ID>IN_0</ID>636 </input>
<input>
<ID>IN_1</ID>909 </input>
<output>
<ID>OUT</ID>650 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>742</ID>
<type>DE_TO</type>
<position>177,-69.5</position>
<input>
<ID>IN_0</ID>986 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN1</lparam></gate>
<gate>
<ID>381</ID>
<type>AA_AND2</type>
<position>197.5,-120.5</position>
<input>
<ID>IN_0</ID>642 </input>
<input>
<ID>IN_1</ID>643 </input>
<output>
<ID>OUT</ID>655 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>382</ID>
<type>AA_AND2</type>
<position>197.5,-126.5</position>
<input>
<ID>IN_0</ID>645 </input>
<input>
<ID>IN_1</ID>913 </input>
<output>
<ID>OUT</ID>654 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>229</ID>
<type>FF_GND</type>
<position>168,-120</position>
<output>
<ID>OUT_0</ID>504 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>383</ID>
<type>AA_AND2</type>
<position>197.5,-132.5</position>
<input>
<ID>IN_0</ID>647 </input>
<input>
<ID>IN_1</ID>914 </input>
<output>
<ID>OUT</ID>653 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>730</ID>
<type>DA_FROM</type>
<position>192,-200</position>
<input>
<ID>IN_0</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr14</lparam></gate>
<gate>
<ID>384</ID>
<type>DA_FROM</type>
<position>192.5,-93.5</position>
<input>
<ID>IN_0</ID>633 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>689</ID>
<type>DA_FROM</type>
<position>140,-154.5</position>
<input>
<ID>IN_0</ID>934 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr9</lparam></gate>
<gate>
<ID>386</ID>
<type>DA_FROM</type>
<position>192.5,-101.5</position>
<input>
<ID>IN_0</ID>636 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>388</ID>
<type>DA_FROM</type>
<position>192.5,-107.5</position>
<input>
<ID>IN_0</ID>638 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR</lparam></gate>
<gate>
<ID>693</ID>
<type>DA_FROM</type>
<position>140,-178.5</position>
<input>
<ID>IN_0</ID>938 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac8</lparam></gate>
<gate>
<ID>390</ID>
<type>DA_FROM</type>
<position>192.5,-113.5</position>
<input>
<ID>IN_0</ID>640 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>392</ID>
<type>DA_FROM</type>
<position>192.5,-119.5</position>
<input>
<ID>IN_0</ID>642 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>394</ID>
<type>AE_SMALL_INVERTER</type>
<position>192.5,-121.5</position>
<input>
<ID>IN_0</ID>912 </input>
<output>
<ID>OUT_0</ID>643 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>559</ID>
<type>AA_AND2</type>
<position>197,-199</position>
<input>
<ID>IN_0</ID>830 </input>
<input>
<ID>IN_1</ID>974 </input>
<output>
<ID>OUT</ID>843 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>395</ID>
<type>DA_FROM</type>
<position>192.5,-125.5</position>
<input>
<ID>IN_0</ID>645 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>397</ID>
<type>DA_FROM</type>
<position>192.5,-131.5</position>
<input>
<ID>IN_0</ID>647 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>732</ID>
<type>DA_FROM</type>
<position>188,-212</position>
<input>
<ID>IN_0</ID>976 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac14</lparam></gate>
<gate>
<ID>547</ID>
<type>DA_FROM</type>
<position>88.5,-210</position>
<input>
<ID>IN_0</ID>786 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>399</ID>
<type>DE_OR8</type>
<position>223,-115</position>
<input>
<ID>IN_0</ID>649 </input>
<input>
<ID>IN_1</ID>650 </input>
<input>
<ID>IN_2</ID>651 </input>
<input>
<ID>IN_3</ID>652 </input>
<input>
<ID>IN_4</ID>500 </input>
<input>
<ID>IN_5</ID>653 </input>
<input>
<ID>IN_6</ID>654 </input>
<input>
<ID>IN_7</ID>655 </input>
<output>
<ID>OUT</ID>991 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>577</ID>
<type>AE_SMALL_INVERTER</type>
<position>140,-212</position>
<input>
<ID>IN_0</ID>968 </input>
<output>
<ID>OUT_0</ID>811 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>401</ID>
<type>AA_AND3</type>
<position>249,-95.5</position>
<input>
<ID>IN_0</ID>657 </input>
<input>
<ID>IN_1</ID>915 </input>
<input>
<ID>IN_2</ID>916 </input>
<output>
<ID>OUT</ID>673 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>736</ID>
<type>DA_FROM</type>
<position>243.5,-188</position>
<input>
<ID>IN_0</ID>980 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac15</lparam></gate>
<gate>
<ID>402</ID>
<type>AA_AND2</type>
<position>249,-102.5</position>
<input>
<ID>IN_0</ID>660 </input>
<input>
<ID>IN_1</ID>917 </input>
<output>
<ID>OUT</ID>674 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>403</ID>
<type>AA_AND2</type>
<position>249,-108.5</position>
<input>
<ID>IN_0</ID>662 </input>
<input>
<ID>IN_1</ID>918 </input>
<output>
<ID>OUT</ID>675 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>404</ID>
<type>AA_AND2</type>
<position>249,-114.5</position>
<input>
<ID>IN_0</ID>664 </input>
<input>
<ID>IN_1</ID>919 </input>
<output>
<ID>OUT</ID>676 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>405</ID>
<type>DA_FROM</type>
<position>244,-131.5</position>
<input>
<ID>IN_0</ID>671 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>740</ID>
<type>DA_FROM</type>
<position>239.5,-212</position>
<input>
<ID>IN_0</ID>984 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac15</lparam></gate>
<gate>
<ID>406</ID>
<type>AA_AND2</type>
<position>249,-120.5</position>
<input>
<ID>IN_0</ID>666 </input>
<input>
<ID>IN_1</ID>667 </input>
<output>
<ID>OUT</ID>679 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>407</ID>
<type>AA_AND2</type>
<position>249,-126.5</position>
<input>
<ID>IN_0</ID>669 </input>
<input>
<ID>IN_1</ID>921 </input>
<output>
<ID>OUT</ID>678 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>408</ID>
<type>AA_AND2</type>
<position>249,-132.5</position>
<input>
<ID>IN_0</ID>671 </input>
<input>
<ID>IN_1</ID>922 </input>
<output>
<ID>OUT</ID>677 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>585</ID>
<type>AA_AND2</type>
<position>197,-217</position>
<input>
<ID>IN_0</ID>837 </input>
<input>
<ID>IN_1</ID>977 </input>
<output>
<ID>OUT</ID>846 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>409</ID>
<type>DA_FROM</type>
<position>244,-93.5</position>
<input>
<ID>IN_0</ID>657 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>744</ID>
<type>DE_TO</type>
<position>280.5,-69.5</position>
<input>
<ID>IN_0</ID>988 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN3</lparam></gate>
<gate>
<ID>575</ID>
<type>DA_FROM</type>
<position>140,-210</position>
<input>
<ID>IN_0</ID>810 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>412</ID>
<type>DA_FROM</type>
<position>244,-101.5</position>
<input>
<ID>IN_0</ID>660 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>589</ID>
<type>DA_FROM</type>
<position>192,-192</position>
<input>
<ID>IN_0</ID>828 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>414</ID>
<type>DA_FROM</type>
<position>244,-107.5</position>
<input>
<ID>IN_0</ID>662 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR</lparam></gate>
<gate>
<ID>563</ID>
<type>AA_AND2</type>
<position>145,-211</position>
<input>
<ID>IN_0</ID>810 </input>
<input>
<ID>IN_1</ID>811 </input>
<output>
<ID>OUT</ID>823 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>416</ID>
<type>DA_FROM</type>
<position>244,-113.5</position>
<input>
<ID>IN_0</ID>664 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>593</ID>
<type>DA_FROM</type>
<position>192,-210</position>
<input>
<ID>IN_0</ID>834 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>418</ID>
<type>DA_FROM</type>
<position>244,-119.5</position>
<input>
<ID>IN_0</ID>666 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>420</ID>
<type>AE_SMALL_INVERTER</type>
<position>244,-121.5</position>
<input>
<ID>IN_0</ID>920 </input>
<output>
<ID>OUT_0</ID>667 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>421</ID>
<type>DA_FROM</type>
<position>244,-125.5</position>
<input>
<ID>IN_0</ID>669 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>756</ID>
<type>DE_TO</type>
<position>280,-205.5</position>
<input>
<ID>IN_0</ID>1000 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN15</lparam></gate>
<gate>
<ID>571</ID>
<type>DA_FROM</type>
<position>140,-198</position>
<input>
<ID>IN_0</ID>806 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR</lparam></gate>
<gate>
<ID>424</ID>
<type>DE_OR8</type>
<position>274.5,-115</position>
<input>
<ID>IN_0</ID>673 </input>
<input>
<ID>IN_1</ID>674 </input>
<input>
<ID>IN_2</ID>675 </input>
<input>
<ID>IN_3</ID>676 </input>
<input>
<ID>IN_4</ID>486 </input>
<input>
<ID>IN_5</ID>677 </input>
<input>
<ID>IN_6</ID>678 </input>
<input>
<ID>IN_7</ID>679 </input>
<output>
<ID>OUT</ID>992 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>428</ID>
<type>AA_AND2</type>
<position>197,-205</position>
<input>
<ID>IN_0</ID>832 </input>
<input>
<ID>IN_1</ID>975 </input>
<output>
<ID>OUT</ID>844 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>605</ID>
<type>AA_AND2</type>
<position>248.5,-205</position>
<input>
<ID>IN_0</ID>856 </input>
<input>
<ID>IN_1</ID>983 </input>
<output>
<ID>OUT</ID>868 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>430</ID>
<type>AA_AND3</type>
<position>93.5,-140.5</position>
<input>
<ID>IN_0</ID>681 </input>
<input>
<ID>IN_1</ID>923 </input>
<input>
<ID>IN_2</ID>924 </input>
<output>
<ID>OUT</ID>697 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>432</ID>
<type>AA_AND2</type>
<position>93.5,-147.5</position>
<input>
<ID>IN_0</ID>684 </input>
<input>
<ID>IN_1</ID>925 </input>
<output>
<ID>OUT</ID>698 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>609</ID>
<type>AA_AND2</type>
<position>248.5,-223</position>
<input>
<ID>IN_0</ID>863 </input>
<input>
<ID>IN_1</ID>985 </input>
<output>
<ID>OUT</ID>869 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>433</ID>
<type>AA_AND2</type>
<position>93.5,-153.5</position>
<input>
<ID>IN_0</ID>686 </input>
<input>
<ID>IN_1</ID>926 </input>
<output>
<ID>OUT</ID>699 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>640</ID>
<type>DA_FROM</type>
<position>244,-70</position>
<input>
<ID>IN_0</ID>887 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr3</lparam></gate>
<gate>
<ID>434</ID>
<type>AA_AND2</type>
<position>93.5,-159.5</position>
<input>
<ID>IN_0</ID>688 </input>
<input>
<ID>IN_1</ID>927 </input>
<output>
<ID>OUT</ID>700 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>435</ID>
<type>AA_AND2</type>
<position>93.5,-165.5</position>
<input>
<ID>IN_0</ID>690 </input>
<input>
<ID>IN_1</ID>691 </input>
<output>
<ID>OUT</ID>703 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>436</ID>
<type>AA_AND2</type>
<position>93.5,-171.5</position>
<input>
<ID>IN_0</ID>693 </input>
<input>
<ID>IN_1</ID>929 </input>
<output>
<ID>OUT</ID>702 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>613</ID>
<type>DA_FROM</type>
<position>243.5,-192</position>
<input>
<ID>IN_0</ID>852 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>437</ID>
<type>AA_AND2</type>
<position>93.5,-177.5</position>
<input>
<ID>IN_0</ID>695 </input>
<input>
<ID>IN_1</ID>930 </input>
<output>
<ID>OUT</ID>701 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>644</ID>
<type>DA_FROM</type>
<position>89,-95.5</position>
<input>
<ID>IN_0</ID>891 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr4</lparam></gate>
<gate>
<ID>438</ID>
<type>DA_FROM</type>
<position>88.5,-138.5</position>
<input>
<ID>IN_0</ID>681 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>441</ID>
<type>DA_FROM</type>
<position>88.5,-146.5</position>
<input>
<ID>IN_0</ID>684 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>648</ID>
<type>DA_FROM</type>
<position>89,-115.5</position>
<input>
<ID>IN_0</ID>895 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr4</lparam></gate>
<gate>
<ID>443</ID>
<type>DA_FROM</type>
<position>88.5,-152.5</position>
<input>
<ID>IN_0</ID>686 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR</lparam></gate>
<gate>
<ID>621</ID>
<type>DA_FROM</type>
<position>243.5,-216</position>
<input>
<ID>IN_0</ID>861 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>445</ID>
<type>DA_FROM</type>
<position>88.5,-158.5</position>
<input>
<ID>IN_0</ID>688 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>652</ID>
<type>DA_FROM</type>
<position>140.5,-95.5</position>
<input>
<ID>IN_0</ID>899 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr5</lparam></gate>
<gate>
<ID>447</ID>
<type>DA_FROM</type>
<position>88.5,-164.5</position>
<input>
<ID>IN_0</ID>690 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>449</ID>
<type>AE_SMALL_INVERTER</type>
<position>88.5,-166.5</position>
<input>
<ID>IN_0</ID>928 </input>
<output>
<ID>OUT_0</ID>691 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>450</ID>
<type>DA_FROM</type>
<position>88.5,-170.5</position>
<input>
<ID>IN_0</ID>693 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>452</ID>
<type>DA_FROM</type>
<position>88.5,-176.5</position>
<input>
<ID>IN_0</ID>695 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>454</ID>
<type>DE_OR8</type>
<position>119,-160</position>
<input>
<ID>IN_0</ID>697 </input>
<input>
<ID>IN_1</ID>698 </input>
<input>
<ID>IN_2</ID>699 </input>
<input>
<ID>IN_3</ID>700 </input>
<input>
<ID>IN_4</ID>328 </input>
<input>
<ID>IN_5</ID>701 </input>
<input>
<ID>IN_6</ID>702 </input>
<input>
<ID>IN_7</ID>703 </input>
<output>
<ID>OUT</ID>993 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>603</ID>
<type>AA_AND2</type>
<position>248.5,-193</position>
<input>
<ID>IN_0</ID>852 </input>
<input>
<ID>IN_1</ID>981 </input>
<output>
<ID>OUT</ID>866 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>457</ID>
<type>AA_AND3</type>
<position>145,-140.5</position>
<input>
<ID>IN_0</ID>705 </input>
<input>
<ID>IN_1</ID>931 </input>
<input>
<ID>IN_2</ID>932 </input>
<output>
<ID>OUT</ID>721 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>458</ID>
<type>AA_AND2</type>
<position>145,-147.5</position>
<input>
<ID>IN_0</ID>708 </input>
<input>
<ID>IN_1</ID>933 </input>
<output>
<ID>OUT</ID>722 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>460</ID>
<type>AA_AND2</type>
<position>145,-153.5</position>
<input>
<ID>IN_0</ID>710 </input>
<input>
<ID>IN_1</ID>934 </input>
<output>
<ID>OUT</ID>723 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>461</ID>
<type>AA_AND2</type>
<position>145,-159.5</position>
<input>
<ID>IN_0</ID>712 </input>
<input>
<ID>IN_1</ID>935 </input>
<output>
<ID>OUT</ID>724 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>462</ID>
<type>DA_FROM</type>
<position>140,-176.5</position>
<input>
<ID>IN_0</ID>719 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>463</ID>
<type>AA_AND2</type>
<position>145,-165.5</position>
<input>
<ID>IN_0</ID>714 </input>
<input>
<ID>IN_1</ID>715 </input>
<output>
<ID>OUT</ID>727 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>464</ID>
<type>AA_AND2</type>
<position>145,-171.5</position>
<input>
<ID>IN_0</ID>717 </input>
<input>
<ID>IN_1</ID>937 </input>
<output>
<ID>OUT</ID>726 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>641</ID>
<type>DA_FROM</type>
<position>240,-76</position>
<input>
<ID>IN_0</ID>888 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac3</lparam></gate>
<gate>
<ID>466</ID>
<type>DA_FROM</type>
<position>140,-138.5</position>
<input>
<ID>IN_0</ID>705 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>631</ID>
<type>DA_FROM</type>
<position>192.5,-70</position>
<input>
<ID>IN_0</ID>878 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr2</lparam></gate>
<gate>
<ID>645</ID>
<type>DA_FROM</type>
<position>89,-97.5</position>
<input>
<ID>IN_0</ID>892 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac4</lparam></gate>
<gate>
<ID>649</ID>
<type>DA_FROM</type>
<position>85,-121.5</position>
<input>
<ID>IN_0</ID>896 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac4</lparam></gate>
<gate>
<ID>474</ID>
<type>DE_TO</type>
<position>117.5,-24</position>
<input>
<ID>IN_0</ID>608 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr12</lparam></gate>
<gate>
<ID>639</ID>
<type>DA_FROM</type>
<position>244,-64</position>
<input>
<ID>IN_0</ID>886 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr3</lparam></gate>
<gate>
<ID>653</ID>
<type>DA_FROM</type>
<position>140.5,-97.5</position>
<input>
<ID>IN_0</ID>900 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac5</lparam></gate>
<gate>
<ID>478</ID>
<type>DA_FROM</type>
<position>140,-170.5</position>
<input>
<ID>IN_0</ID>717 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>627</ID>
<type>DA_FROM</type>
<position>192.5,-50</position>
<input>
<ID>IN_0</ID>874 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr2</lparam></gate>
<gate>
<ID>657</ID>
<type>DA_FROM</type>
<position>136.5,-121.5</position>
<input>
<ID>IN_0</ID>904 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac5</lparam></gate>
<gate>
<ID>482</ID>
<type>DE_TO</type>
<position>117.5,-28</position>
<input>
<ID>IN_0</ID>608 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr14</lparam></gate>
<gate>
<ID>519</ID>
<type>DA_FROM</type>
<position>243.5,-152.5</position>
<input>
<ID>IN_0</ID>758 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR</lparam></gate>
<gate>
<ID>483</ID>
<type>AA_AND3</type>
<position>197,-140.5</position>
<input>
<ID>IN_0</ID>729 </input>
<input>
<ID>IN_1</ID>939 </input>
<input>
<ID>IN_2</ID>940 </input>
<output>
<ID>OUT</ID>745 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>484</ID>
<type>AA_AND2</type>
<position>197,-147.5</position>
<input>
<ID>IN_0</ID>732 </input>
<input>
<ID>IN_1</ID>941 </input>
<output>
<ID>OUT</ID>746 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>661</ID>
<type>DA_FROM</type>
<position>192.5,-97.5</position>
<input>
<ID>IN_0</ID>908 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac6</lparam></gate>
<gate>
<ID>486</ID>
<type>AA_AND2</type>
<position>197,-165.5</position>
<input>
<ID>IN_0</ID>738 </input>
<input>
<ID>IN_1</ID>739 </input>
<output>
<ID>OUT</ID>751 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>635</ID>
<type>DA_FROM</type>
<position>192.5,-88</position>
<input>
<ID>IN_0</ID>882 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac1</lparam></gate>
<gate>
<ID>488</ID>
<type>AA_AND2</type>
<position>197,-177.5</position>
<input>
<ID>IN_0</ID>743 </input>
<input>
<ID>IN_1</ID>946 </input>
<output>
<ID>OUT</ID>749 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>665</ID>
<type>DA_FROM</type>
<position>188.5,-121.5</position>
<input>
<ID>IN_0</ID>912 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac6</lparam></gate>
<gate>
<ID>489</ID>
<type>DA_FROM</type>
<position>192,-138.5</position>
<input>
<ID>IN_0</ID>729 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>491</ID>
<type>DA_FROM</type>
<position>192,-146.5</position>
<input>
<ID>IN_0</ID>732 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>492</ID>
<type>DE_TO</type>
<position>117.5,-30</position>
<input>
<ID>IN_0</ID>608 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr15</lparam></gate>
<gate>
<ID>669</ID>
<type>DA_FROM</type>
<position>244,-97.5</position>
<input>
<ID>IN_0</ID>916 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac7</lparam></gate>
<gate>
<ID>493</ID>
<type>DA_FROM</type>
<position>192,-152.5</position>
<input>
<ID>IN_0</ID>734 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR</lparam></gate>
<gate>
<ID>495</ID>
<type>DA_FROM</type>
<position>192,-158.5</position>
<input>
<ID>IN_0</ID>736 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>673</ID>
<type>DA_FROM</type>
<position>240,-121.5</position>
<input>
<ID>IN_0</ID>920 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac7</lparam></gate>
<gate>
<ID>497</ID>
<type>DA_FROM</type>
<position>192,-164.5</position>
<input>
<ID>IN_0</ID>738 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>704</ID>
<type>DA_FROM</type>
<position>243.5,-142.5</position>
<input>
<ID>IN_0</ID>948 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac11</lparam></gate>
<gate>
<ID>535</ID>
<type>AA_AND2</type>
<position>93.5,-211</position>
<input>
<ID>IN_0</ID>786 </input>
<input>
<ID>IN_1</ID>787 </input>
<output>
<ID>OUT</ID>799 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>500</ID>
<type>DA_FROM</type>
<position>192,-170.5</position>
<input>
<ID>IN_0</ID>741 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>677</ID>
<type>DA_FROM</type>
<position>88.5,-142.5</position>
<input>
<ID>IN_0</ID>924 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac8</lparam></gate>
<gate>
<ID>502</ID>
<type>DA_FROM</type>
<position>192,-176.5</position>
<input>
<ID>IN_0</ID>743 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>523</ID>
<type>DA_FROM</type>
<position>243.5,-164.5</position>
<input>
<ID>IN_0</ID>762 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>504</ID>
<type>DE_OR8</type>
<position>222.5,-160</position>
<input>
<ID>IN_0</ID>745 </input>
<input>
<ID>IN_1</ID>746 </input>
<input>
<ID>IN_2</ID>747 </input>
<input>
<ID>IN_3</ID>748 </input>
<input>
<ID>IN_4</ID>471 </input>
<input>
<ID>IN_5</ID>749 </input>
<input>
<ID>IN_6</ID>750 </input>
<input>
<ID>IN_7</ID>751 </input>
<output>
<ID>OUT</ID>995 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>681</ID>
<type>DA_FROM</type>
<position>84.5,-166.5</position>
<input>
<ID>IN_0</ID>928 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac8</lparam></gate>
<gate>
<ID>712</ID>
<type>DA_FROM</type>
<position>88.5,-188</position>
<input>
<ID>IN_0</ID>956 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac12</lparam></gate>
<gate>
<ID>506</ID>
<type>AA_AND3</type>
<position>248.5,-140.5</position>
<input>
<ID>IN_0</ID>753 </input>
<input>
<ID>IN_1</ID>947 </input>
<input>
<ID>IN_2</ID>948 </input>
<output>
<ID>OUT</ID>769 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>543</ID>
<type>DA_FROM</type>
<position>88.5,-198</position>
<input>
<ID>IN_0</ID>782 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR</lparam></gate>
<gate>
<ID>507</ID>
<type>AA_AND2</type>
<position>248.5,-147.5</position>
<input>
<ID>IN_0</ID>756 </input>
<input>
<ID>IN_1</ID>949 </input>
<output>
<ID>OUT</ID>770 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>508</ID>
<type>AA_AND2</type>
<position>248.5,-153.5</position>
<input>
<ID>IN_0</ID>758 </input>
<input>
<ID>IN_1</ID>950 </input>
<output>
<ID>OUT</ID>771 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>509</ID>
<type>AA_AND2</type>
<position>248.5,-159.5</position>
<input>
<ID>IN_0</ID>760 </input>
<input>
<ID>IN_1</ID>951 </input>
<output>
<ID>OUT</ID>772 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>716</ID>
<type>DA_FROM</type>
<position>84.5,-212</position>
<input>
<ID>IN_0</ID>960 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac12</lparam></gate>
<gate>
<ID>510</ID>
<type>DA_FROM</type>
<position>243.5,-176.5</position>
<input>
<ID>IN_0</ID>767 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>531</ID>
<type>AA_AND3</type>
<position>93.5,-186</position>
<input>
<ID>IN_0</ID>777 </input>
<input>
<ID>IN_1</ID>955 </input>
<input>
<ID>IN_2</ID>956 </input>
<output>
<ID>OUT</ID>793 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>514</ID>
<type>DA_FROM</type>
<position>243.5,-138.5</position>
<input>
<ID>IN_0</ID>753 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>526</ID>
<type>DA_FROM</type>
<position>243.5,-170.5</position>
<input>
<ID>IN_0</ID>765 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>532</ID>
<type>AA_AND2</type>
<position>93.5,-193</position>
<input>
<ID>IN_0</ID>780 </input>
<input>
<ID>IN_1</ID>957 </input>
<output>
<ID>OUT</ID>794 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>534</ID>
<type>AA_AND2</type>
<position>93.5,-205</position>
<input>
<ID>IN_0</ID>784 </input>
<input>
<ID>IN_1</ID>959 </input>
<output>
<ID>OUT</ID>796 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>536</ID>
<type>AA_AND2</type>
<position>93.5,-217</position>
<input>
<ID>IN_0</ID>789 </input>
<input>
<ID>IN_1</ID>961 </input>
<output>
<ID>OUT</ID>798 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>538</ID>
<type>DA_FROM</type>
<position>88.5,-184</position>
<input>
<ID>IN_0</ID>777 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>552</ID>
<type>DA_FROM</type>
<position>88.5,-222</position>
<input>
<ID>IN_0</ID>791 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>554</ID>
<type>DE_OR8</type>
<position>119,-205.5</position>
<input>
<ID>IN_0</ID>793 </input>
<input>
<ID>IN_1</ID>794 </input>
<input>
<ID>IN_2</ID>795 </input>
<input>
<ID>IN_3</ID>796 </input>
<input>
<ID>IN_4</ID>323 </input>
<input>
<ID>IN_5</ID>797 </input>
<input>
<ID>IN_6</ID>798 </input>
<input>
<ID>IN_7</ID>799 </input>
<output>
<ID>OUT</ID>997 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>224</ID>
<type>FF_GND</type>
<position>271,-165</position>
<output>
<ID>OUT_0</ID>472 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>560</ID>
<type>AA_AND2</type>
<position>145,-199</position>
<input>
<ID>IN_0</ID>806 </input>
<input>
<ID>IN_1</ID>966 </input>
<output>
<ID>OUT</ID>819 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>564</ID>
<type>AA_AND2</type>
<position>145,-217</position>
<input>
<ID>IN_0</ID>813 </input>
<input>
<ID>IN_1</ID>969 </input>
<output>
<ID>OUT</ID>822 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>578</ID>
<type>DA_FROM</type>
<position>140,-216</position>
<input>
<ID>IN_0</ID>813 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>582</ID>
<type>AA_AND3</type>
<position>197,-186</position>
<input>
<ID>IN_0</ID>825 </input>
<input>
<ID>IN_1</ID>971 </input>
<input>
<ID>IN_2</ID>972 </input>
<output>
<ID>OUT</ID>841 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>583</ID>
<type>AA_AND2</type>
<position>197,-193</position>
<input>
<ID>IN_0</ID>828 </input>
<input>
<ID>IN_1</ID>973 </input>
<output>
<ID>OUT</ID>842 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>586</ID>
<type>AA_AND2</type>
<position>197,-223</position>
<input>
<ID>IN_0</ID>839 </input>
<input>
<ID>IN_1</ID>978 </input>
<output>
<ID>OUT</ID>845 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>587</ID>
<type>DA_FROM</type>
<position>192,-184</position>
<input>
<ID>IN_0</ID>825 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>590</ID>
<type>DA_FROM</type>
<position>192,-198</position>
<input>
<ID>IN_0</ID>830 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR</lparam></gate>
<gate>
<ID>595</ID>
<type>AE_SMALL_INVERTER</type>
<position>192,-212</position>
<input>
<ID>IN_0</ID>976 </input>
<output>
<ID>OUT_0</ID>835 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>598</ID>
<type>DA_FROM</type>
<position>192,-222</position>
<input>
<ID>IN_0</ID>839 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>602</ID>
<type>AA_AND3</type>
<position>248.5,-186</position>
<input>
<ID>IN_0</ID>849 </input>
<input>
<ID>IN_1</ID>979 </input>
<input>
<ID>IN_2</ID>980 </input>
<output>
<ID>OUT</ID>865 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>606</ID>
<type>DA_FROM</type>
<position>243.5,-222</position>
<input>
<ID>IN_0</ID>863 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>607</ID>
<type>AA_AND2</type>
<position>248.5,-211</position>
<input>
<ID>IN_0</ID>858 </input>
<input>
<ID>IN_1</ID>859 </input>
<output>
<ID>OUT</ID>871 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>610</ID>
<type>DA_FROM</type>
<position>243.5,-184</position>
<input>
<ID>IN_0</ID>849 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>614</ID>
<type>DA_FROM</type>
<position>243.5,-198</position>
<input>
<ID>IN_0</ID>854 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR</lparam></gate>
<gate>
<ID>618</ID>
<type>DA_FROM</type>
<position>243.5,-210</position>
<input>
<ID>IN_0</ID>858 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>622</ID>
<type>DA_FROM</type>
<position>243.5,-218</position>
<input>
<ID>IN_0</ID>862 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac0</lparam></gate>
<gate>
<ID>630</ID>
<type>DA_FROM</type>
<position>192.5,-64</position>
<input>
<ID>IN_0</ID>877 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr2</lparam></gate>
<gate>
<ID>634</ID>
<type>DA_FROM</type>
<position>140.5,-88</position>
<input>
<ID>IN_0</ID>881 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac0</lparam></gate>
<gate>
<ID>638</ID>
<type>DA_FROM</type>
<position>244,-58</position>
<input>
<ID>IN_0</ID>885 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add3</lparam></gate>
<gate>
<ID>643</ID>
<type>DA_FROM</type>
<position>244,-88</position>
<input>
<ID>IN_0</ID>890 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac2</lparam></gate>
<gate>
<ID>647</ID>
<type>DA_FROM</type>
<position>89,-109.5</position>
<input>
<ID>IN_0</ID>894 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr4</lparam></gate>
<gate>
<ID>651</ID>
<type>DA_FROM</type>
<position>89,-133.5</position>
<input>
<ID>IN_0</ID>898 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac3</lparam></gate>
<gate>
<ID>654</ID>
<type>DA_FROM</type>
<position>140.5,-103.5</position>
<input>
<ID>IN_0</ID>901 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add5</lparam></gate>
<gate>
<ID>655</ID>
<type>DA_FROM</type>
<position>140.5,-109.5</position>
<input>
<ID>IN_0</ID>902 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr5</lparam></gate>
<gate>
<ID>658</ID>
<type>DA_FROM</type>
<position>140.5,-127.5</position>
<input>
<ID>IN_0</ID>905 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac6</lparam></gate>
<gate>
<ID>659</ID>
<type>DA_FROM</type>
<position>140.5,-133.5</position>
<input>
<ID>IN_0</ID>906 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac4</lparam></gate>
<gate>
<ID>663</ID>
<type>DA_FROM</type>
<position>192.5,-109.5</position>
<input>
<ID>IN_0</ID>910 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr6</lparam></gate>
<gate>
<ID>666</ID>
<type>DA_FROM</type>
<position>192.5,-127.5</position>
<input>
<ID>IN_0</ID>913 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac7</lparam></gate>
<gate>
<ID>667</ID>
<type>DA_FROM</type>
<position>192.5,-133.5</position>
<input>
<ID>IN_0</ID>914 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac5</lparam></gate>
<gate>
<ID>671</ID>
<type>DA_FROM</type>
<position>244,-109.5</position>
<input>
<ID>IN_0</ID>918 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr7</lparam></gate>
<gate>
<ID>672</ID>
<type>DA_FROM</type>
<position>244,-115.5</position>
<input>
<ID>IN_0</ID>919 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr7</lparam></gate>
<gate>
<ID>674</ID>
<type>DA_FROM</type>
<position>244,-127.5</position>
<input>
<ID>IN_0</ID>921 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac8</lparam></gate>
<gate>
<ID>675</ID>
<type>DA_FROM</type>
<position>244,-133.5</position>
<input>
<ID>IN_0</ID>922 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac6</lparam></gate>
<gate>
<ID>676</ID>
<type>DA_FROM</type>
<position>88.5,-140.5</position>
<input>
<ID>IN_0</ID>923 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr8</lparam></gate>
<gate>
<ID>678</ID>
<type>DA_FROM</type>
<position>88.5,-148.5</position>
<input>
<ID>IN_0</ID>925 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add8</lparam></gate>
<gate>
<ID>679</ID>
<type>DA_FROM</type>
<position>88.5,-154.5</position>
<input>
<ID>IN_0</ID>926 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr8</lparam></gate>
<gate>
<ID>682</ID>
<type>DA_FROM</type>
<position>88.5,-172.5</position>
<input>
<ID>IN_0</ID>929 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac9</lparam></gate>
<gate>
<ID>683</ID>
<type>DA_FROM</type>
<position>88.5,-178.5</position>
<input>
<ID>IN_0</ID>930 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac7</lparam></gate>
<gate>
<ID>686</ID>
<type>DA_FROM</type>
<position>140,-140.5</position>
<input>
<ID>IN_0</ID>931 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr9</lparam></gate>
<gate>
<ID>687</ID>
<type>DA_FROM</type>
<position>140,-142.5</position>
<input>
<ID>IN_0</ID>932 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac9</lparam></gate>
<gate>
<ID>690</ID>
<type>DA_FROM</type>
<position>140,-160.5</position>
<input>
<ID>IN_0</ID>935 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr9</lparam></gate>
<gate>
<ID>691</ID>
<type>DA_FROM</type>
<position>136,-166.5</position>
<input>
<ID>IN_0</ID>936 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac9</lparam></gate>
<gate>
<ID>694</ID>
<type>DA_FROM</type>
<position>192,-140.5</position>
<input>
<ID>IN_0</ID>939 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr10</lparam></gate>
<gate>
<ID>695</ID>
<type>DA_FROM</type>
<position>192,-142.5</position>
<input>
<ID>IN_0</ID>940 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac10</lparam></gate>
<gate>
<ID>698</ID>
<type>DA_FROM</type>
<position>192,-154.5</position>
<input>
<ID>IN_0</ID>942 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr10</lparam></gate>
<gate>
<ID>699</ID>
<type>DA_FROM</type>
<position>192,-160.5</position>
<input>
<ID>IN_0</ID>943 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr10</lparam></gate>
<gate>
<ID>700</ID>
<type>DA_FROM</type>
<position>188,-166.5</position>
<input>
<ID>IN_0</ID>944 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac10</lparam></gate>
<gate>
<ID>701</ID>
<type>DA_FROM</type>
<position>192,-172.5</position>
<input>
<ID>IN_0</ID>945 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac11</lparam></gate>
<gate>
<ID>702</ID>
<type>DA_FROM</type>
<position>192,-178.5</position>
<input>
<ID>IN_0</ID>946 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac9</lparam></gate>
<gate>
<ID>703</ID>
<type>DA_FROM</type>
<position>243.5,-140.5</position>
<input>
<ID>IN_0</ID>947 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr11</lparam></gate>
<gate>
<ID>705</ID>
<type>DA_FROM</type>
<position>243.5,-148.5</position>
<input>
<ID>IN_0</ID>949 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add11</lparam></gate>
<gate>
<ID>707</ID>
<type>DA_FROM</type>
<position>243.5,-160.5</position>
<input>
<ID>IN_0</ID>951 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr11</lparam></gate>
<gate>
<ID>708</ID>
<type>DA_FROM</type>
<position>239.5,-166.5</position>
<input>
<ID>IN_0</ID>952 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac11</lparam></gate>
<gate>
<ID>709</ID>
<type>DA_FROM</type>
<position>243.5,-172.5</position>
<input>
<ID>IN_0</ID>953 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac12</lparam></gate>
<gate>
<ID>713</ID>
<type>DA_FROM</type>
<position>88.5,-194</position>
<input>
<ID>IN_0</ID>957 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add12</lparam></gate>
<gate>
<ID>714</ID>
<type>DA_FROM</type>
<position>88.5,-200</position>
<input>
<ID>IN_0</ID>958 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr12</lparam></gate>
<gate>
<ID>715</ID>
<type>DA_FROM</type>
<position>88.5,-206</position>
<input>
<ID>IN_0</ID>959 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr12</lparam></gate>
<gate>
<ID>717</ID>
<type>DA_FROM</type>
<position>88.5,-218</position>
<input>
<ID>IN_0</ID>961 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac13</lparam></gate>
<gate>
<ID>719</ID>
<type>DA_FROM</type>
<position>140,-186</position>
<input>
<ID>IN_0</ID>963 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr13</lparam></gate>
<gate>
<ID>720</ID>
<type>DA_FROM</type>
<position>140,-188</position>
<input>
<ID>IN_0</ID>964 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac13</lparam></gate>
<gate>
<ID>721</ID>
<type>DA_FROM</type>
<position>140,-194</position>
<input>
<ID>IN_0</ID>965 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add13</lparam></gate>
<gate>
<ID>722</ID>
<type>DA_FROM</type>
<position>140,-200</position>
<input>
<ID>IN_0</ID>966 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr13</lparam></gate>
<gate>
<ID>724</ID>
<type>DA_FROM</type>
<position>136,-212</position>
<input>
<ID>IN_0</ID>968 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac13</lparam></gate>
<gate>
<ID>725</ID>
<type>DA_FROM</type>
<position>140,-218</position>
<input>
<ID>IN_0</ID>969 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac14</lparam></gate>
<gate>
<ID>726</ID>
<type>DA_FROM</type>
<position>140,-224</position>
<input>
<ID>IN_0</ID>970 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac12</lparam></gate>
<gate>
<ID>727</ID>
<type>DA_FROM</type>
<position>192,-186</position>
<input>
<ID>IN_0</ID>971 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr14</lparam></gate>
<gate>
<ID>728</ID>
<type>DA_FROM</type>
<position>192,-188</position>
<input>
<ID>IN_0</ID>972 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac14</lparam></gate>
<gate>
<ID>729</ID>
<type>DA_FROM</type>
<position>192,-194</position>
<input>
<ID>IN_0</ID>973 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add14</lparam></gate>
<gate>
<ID>733</ID>
<type>DA_FROM</type>
<position>192,-218</position>
<input>
<ID>IN_0</ID>977 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac15</lparam></gate>
<gate>
<ID>734</ID>
<type>DA_FROM</type>
<position>192,-224</position>
<input>
<ID>IN_0</ID>978 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac13</lparam></gate>
<gate>
<ID>737</ID>
<type>DA_FROM</type>
<position>243.5,-194</position>
<input>
<ID>IN_0</ID>981 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add15</lparam></gate>
<gate>
<ID>741</ID>
<type>DA_FROM</type>
<position>243.5,-224</position>
<input>
<ID>IN_0</ID>985 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac14</lparam></gate>
<gate>
<ID>745</ID>
<type>DE_TO</type>
<position>125.5,-115</position>
<input>
<ID>IN_0</ID>989 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN4</lparam></gate>
<gate>
<ID>749</ID>
<type>DE_TO</type>
<position>125,-160</position>
<input>
<ID>IN_0</ID>993 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN8</lparam></gate>
<gate>
<ID>752</ID>
<type>DE_TO</type>
<position>280,-160</position>
<input>
<ID>IN_0</ID>996 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN11</lparam></gate>
<gate>
<ID>753</ID>
<type>DE_TO</type>
<position>125,-205.5</position>
<input>
<ID>IN_0</ID>997 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN12</lparam></gate>
<gate>
<ID>755</ID>
<type>DE_TO</type>
<position>228.5,-205.5</position>
<input>
<ID>IN_0</ID>999 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID acIN14</lparam></gate>
<gate>
<ID>144</ID>
<type>FF_GND</type>
<position>271,-210.5</position>
<output>
<ID>OUT_0</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>148</ID>
<type>FF_GND</type>
<position>219.5,-210.5</position>
<output>
<ID>OUT_0</ID>104 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>152</ID>
<type>FF_GND</type>
<position>167.5,-210.5</position>
<output>
<ID>OUT_0</ID>322 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>156</ID>
<type>FF_GND</type>
<position>116,-210.5</position>
<output>
<ID>OUT_0</ID>323 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>164</ID>
<type>FF_GND</type>
<position>116,-165</position>
<output>
<ID>OUT_0</ID>328 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>222</ID>
<type>FF_GND</type>
<position>167.5,-165</position>
<output>
<ID>OUT_0</ID>331 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>442</ID>
<type>DE_TO</type>
<position>117.5,-16</position>
<input>
<ID>IN_0</ID>608 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr8</lparam></gate>
<gate>
<ID>446</ID>
<type>DE_TO</type>
<position>117.5,-18</position>
<input>
<ID>IN_0</ID>608 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr9</lparam></gate>
<gate>
<ID>453</ID>
<type>DE_TO</type>
<position>117.5,-20</position>
<input>
<ID>IN_0</ID>608 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr10</lparam></gate>
<gate>
<ID>456</ID>
<type>DE_TO</type>
<position>117.5,-22</position>
<input>
<ID>IN_0</ID>608 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID inpr11</lparam></gate>
<gate>
<ID>520</ID>
<type>FF_GND</type>
<position>115.5,-32</position>
<output>
<ID>OUT_0</ID>608 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>769 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271,-156.5,271,-140.5</points>
<connection>
<GID>529</GID>
<name>IN_0</name></connection>
<intersection>-140.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>251.5,-140.5,271,-140.5</points>
<connection>
<GID>506</GID>
<name>OUT</name></connection>
<intersection>271 0</intersection></hsegment></shape></wire>
<wire>
<ID>80 </ID>
<shape>
<vsegment>
<ID>3</ID>
<points>57,-24,57,-22</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<connection>
<GID>5</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>889 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-82,246,-82</points>
<connection>
<GID>642</GID>
<name>IN_0</name></connection>
<connection>
<GID>307</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>72 </ID>
<shape>
<vsegment>
<ID>4</ID>
<points>65,-21,65,-19.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<connection>
<GID>5</GID>
<name>OUT_3</name></connection></vsegment></shape></wire>
<wire>
<ID>439 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-53,65,-52.5</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<connection>
<GID>71</GID>
<name>OUT_2</name></connection></vsegment></shape></wire>
<wire>
<ID>971 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-186,194,-186</points>
<connection>
<GID>582</GID>
<name>IN_1</name></connection>
<connection>
<GID>727</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>285 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-26,57,-23</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<connection>
<GID>5</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>516 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-56,142.5,-56</points>
<connection>
<GID>252</GID>
<name>IN_0</name></connection>
<connection>
<GID>261</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>995 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226.5,-160,226.5,-160</points>
<connection>
<GID>751</GID>
<name>IN_0</name></connection>
<connection>
<GID>504</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>78 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-20,57,-20</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<connection>
<GID>37</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>288 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-36,65,-35.5</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<connection>
<GID>49</GID>
<name>OUT_2</name></connection></vsegment></shape></wire>
<wire>
<ID>79 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-22,57,-21</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<connection>
<GID>5</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>988 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278.5,-69.5,278.5,-69.5</points>
<connection>
<GID>324</GID>
<name>OUT</name></connection>
<connection>
<GID>744</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>294 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-37,57,-37</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<connection>
<GID>63</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>796 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96.5,-205,116,-205</points>
<connection>
<GID>534</GID>
<name>OUT</name></connection>
<connection>
<GID>554</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>763 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-166.5,245.5,-166.5</points>
<connection>
<GID>511</GID>
<name>IN_1</name></connection>
<connection>
<GID>525</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>924 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-142.5,90.5,-142.5</points>
<connection>
<GID>430</GID>
<name>IN_2</name></connection>
<connection>
<GID>677</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>77 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-13,57,-11.5</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<connection>
<GID>5</GID>
<name>IN_B_0</name></connection></vsegment></shape></wire>
<wire>
<ID>497 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>102,-22,103.5,-22</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>102 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>102,-22.5,102,-22</points>
<connection>
<GID>138</GID>
<name>OUT_4</name></connection>
<intersection>-22 2</intersection></vsegment></shape></wire>
<wire>
<ID>74 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-14,57,-13.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<connection>
<GID>5</GID>
<name>IN_B_1</name></connection></vsegment></shape></wire>
<wire>
<ID>75 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-15.5,57,-15</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<connection>
<GID>5</GID>
<name>IN_B_2</name></connection></vsegment></shape></wire>
<wire>
<ID>662 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-107.5,246,-107.5</points>
<connection>
<GID>403</GID>
<name>IN_0</name></connection>
<connection>
<GID>414</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>299 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-51.5,65,-51</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<connection>
<GID>71</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>893 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-103.5,91,-103.5</points>
<connection>
<GID>646</GID>
<name>IN_0</name></connection>
<connection>
<GID>327</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>76 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-17.5,57,-16</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<connection>
<GID>5</GID>
<name>IN_B_3</name></connection></vsegment></shape></wire>
<wire>
<ID>608 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-31,115.5,-16</points>
<connection>
<GID>479</GID>
<name>IN_0</name></connection>
<connection>
<GID>474</GID>
<name>IN_0</name></connection>
<connection>
<GID>482</GID>
<name>IN_0</name></connection>
<connection>
<GID>492</GID>
<name>IN_0</name></connection>
<connection>
<GID>442</GID>
<name>IN_0</name></connection>
<connection>
<GID>446</GID>
<name>IN_0</name></connection>
<connection>
<GID>453</GID>
<name>IN_0</name></connection>
<connection>
<GID>456</GID>
<name>IN_0</name></connection>
<connection>
<GID>520</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>975 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-206,194,-206</points>
<connection>
<GID>731</GID>
<name>IN_0</name></connection>
<connection>
<GID>428</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>465 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>60,-10,66,-10</points>
<connection>
<GID>126</GID>
<name>OUT_0</name></connection>
<connection>
<GID>5</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>980 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-188,245.5,-188</points>
<connection>
<GID>736</GID>
<name>IN_0</name></connection>
<connection>
<GID>602</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>286 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-33.5,65,-32</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>916 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-97.5,246,-97.5</points>
<connection>
<GID>401</GID>
<name>IN_2</name></connection>
<connection>
<GID>669</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>69 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-16.5,65,-15</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>636 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-101.5,194.5,-101.5</points>
<connection>
<GID>379</GID>
<name>IN_0</name></connection>
<connection>
<GID>386</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>987 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>227,-69.5,227,-69.5</points>
<connection>
<GID>743</GID>
<name>IN_0</name></connection>
<connection>
<GID>299</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>70 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-17.5,65,-17</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<connection>
<GID>5</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>71 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-19,65,-18.5</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<connection>
<GID>5</GID>
<name>OUT_2</name></connection></vsegment></shape></wire>
<wire>
<ID>955 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-186,90.5,-186</points>
<connection>
<GID>711</GID>
<name>IN_0</name></connection>
<connection>
<GID>531</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>461 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-27,60,-26</points>
<connection>
<GID>49</GID>
<name>carry_in</name></connection>
<connection>
<GID>5</GID>
<name>carry_out</name></connection></vsegment></shape></wire>
<wire>
<ID>440 </ID>
<shape>
<vsegment>
<ID>4</ID>
<points>65,-55,65,-53.5</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<connection>
<GID>71</GID>
<name>OUT_3</name></connection></vsegment></shape></wire>
<wire>
<ID>298 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-50.5,65,-49</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>992 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278.5,-115,278.5,-115</points>
<connection>
<GID>748</GID>
<name>IN_0</name></connection>
<connection>
<GID>424</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>628 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>148.5,-114.5,168,-114.5</points>
<connection>
<GID>356</GID>
<name>OUT</name></connection>
<connection>
<GID>376</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>979 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-186,245.5,-186</points>
<connection>
<GID>735</GID>
<name>IN_0</name></connection>
<connection>
<GID>602</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>293 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-30,57,-28.5</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<connection>
<GID>49</GID>
<name>IN_B_0</name></connection></vsegment></shape></wire>
<wire>
<ID>762 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-164.5,245.5,-164.5</points>
<connection>
<GID>511</GID>
<name>IN_0</name></connection>
<connection>
<GID>523</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>287 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-34.5,65,-34</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<connection>
<GID>49</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>967 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-206,142,-206</points>
<connection>
<GID>723</GID>
<name>IN_0</name></connection>
<connection>
<GID>561</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>457 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-71,57,-71</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<connection>
<GID>112</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>775 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269.5,-165.5,269.5,-160.5</points>
<intersection>-165.5 2</intersection>
<intersection>-160.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>269.5,-160.5,271,-160.5</points>
<connection>
<GID>529</GID>
<name>IN_7</name></connection>
<intersection>269.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>251.5,-165.5,269.5,-165.5</points>
<connection>
<GID>511</GID>
<name>OUT</name></connection>
<intersection>269.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>446 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-56,57,-55</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<connection>
<GID>71</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>97 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271,-209.5,271,-209</points>
<connection>
<GID>624</GID>
<name>IN_4</name></connection>
<connection>
<GID>144</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>944 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190,-166.5,190,-166.5</points>
<connection>
<GID>499</GID>
<name>IN_0</name></connection>
<connection>
<GID>700</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>462 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-44,60,-43</points>
<connection>
<GID>71</GID>
<name>carry_in</name></connection>
<connection>
<GID>49</GID>
<name>carry_out</name></connection></vsegment></shape></wire>
<wire>
<ID>772 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>251.5,-159.5,271,-159.5</points>
<connection>
<GID>509</GID>
<name>OUT</name></connection>
<connection>
<GID>529</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>739 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-166.5,194,-166.5</points>
<connection>
<GID>499</GID>
<name>OUT_0</name></connection>
<connection>
<GID>486</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>623 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-131.5,142.5,-131.5</points>
<connection>
<GID>357</GID>
<name>IN_0</name></connection>
<connection>
<GID>360</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>458 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-73,57,-72</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<connection>
<GID>84</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>797 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-223,115.5,-208</points>
<intersection>-223 2</intersection>
<intersection>-208 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>96.5,-223,115.5,-223</points>
<connection>
<GID>537</GID>
<name>OUT</name></connection>
<intersection>115.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>115.5,-208,116,-208</points>
<connection>
<GID>554</GID>
<name>IN_5</name></connection>
<intersection>115.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>459 </ID>
<shape>
<vsegment>
<ID>3</ID>
<points>57,-75,57,-73</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<connection>
<GID>84</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>765 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-170.5,245.5,-170.5</points>
<connection>
<GID>512</GID>
<name>IN_0</name></connection>
<connection>
<GID>526</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>460 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-77,57,-74</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<connection>
<GID>84</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>786 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-210,90.5,-210</points>
<connection>
<GID>547</GID>
<name>IN_0</name></connection>
<connection>
<GID>535</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>456 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-64,57,-62.5</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<connection>
<GID>84</GID>
<name>IN_B_0</name></connection></vsegment></shape></wire>
<wire>
<ID>453 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-65,57,-64.5</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<connection>
<GID>84</GID>
<name>IN_B_1</name></connection></vsegment></shape></wire>
<wire>
<ID>603 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-113.5,115.5,-108.5</points>
<intersection>-113.5 1</intersection>
<intersection>-108.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115.5,-113.5,116.5,-113.5</points>
<connection>
<GID>349</GID>
<name>IN_2</name></connection>
<intersection>115.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97,-108.5,115.5,-108.5</points>
<connection>
<GID>328</GID>
<name>OUT</name></connection>
<intersection>115.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>454 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-66.5,57,-66</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<connection>
<GID>84</GID>
<name>IN_B_2</name></connection></vsegment></shape></wire>
<wire>
<ID>777 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-184,90.5,-184</points>
<connection>
<GID>531</GID>
<name>IN_0</name></connection>
<connection>
<GID>538</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>455 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-68.5,57,-67</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<connection>
<GID>84</GID>
<name>IN_B_3</name></connection></vsegment></shape></wire>
<wire>
<ID>463 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-61,60,-60</points>
<connection>
<GID>71</GID>
<name>carry_out</name></connection>
<connection>
<GID>84</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>449 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-67.5,65,-66</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>450 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-68.5,65,-68</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<connection>
<GID>84</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>789 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-216,90.5,-216</points>
<connection>
<GID>550</GID>
<name>IN_0</name></connection>
<connection>
<GID>536</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>451 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-70,65,-69.5</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<connection>
<GID>84</GID>
<name>OUT_2</name></connection></vsegment></shape></wire>
<wire>
<ID>782 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-198,90.5,-198</points>
<connection>
<GID>533</GID>
<name>IN_0</name></connection>
<connection>
<GID>543</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>452 </ID>
<shape>
<vsegment>
<ID>4</ID>
<points>65,-72,65,-70.5</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<connection>
<GID>84</GID>
<name>OUT_3</name></connection></vsegment></shape></wire>
<wire>
<ID>794 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-203,115.5,-193</points>
<intersection>-203 1</intersection>
<intersection>-193 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115.5,-203,116,-203</points>
<connection>
<GID>554</GID>
<name>IN_1</name></connection>
<intersection>115.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>96.5,-193,115.5,-193</points>
<connection>
<GID>532</GID>
<name>OUT</name></connection>
<intersection>115.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>464 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-77,60,-77</points>
<connection>
<GID>84</GID>
<name>carry_out</name></connection>
<connection>
<GID>122</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>642 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-119.5,194.5,-119.5</points>
<connection>
<GID>381</GID>
<name>IN_0</name></connection>
<connection>
<GID>392</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>295 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-39,57,-38</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<connection>
<GID>49</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>296 </ID>
<shape>
<vsegment>
<ID>3</ID>
<points>57,-41,57,-39</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<connection>
<GID>49</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>999 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226.5,-205.5,226.5,-205.5</points>
<connection>
<GID>600</GID>
<name>OUT</name></connection>
<connection>
<GID>755</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>297 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-43,57,-40</points>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<connection>
<GID>49</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>920 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242,-121.5,242,-121.5</points>
<connection>
<GID>420</GID>
<name>IN_0</name></connection>
<connection>
<GID>673</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>73 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,-21.5,103,-20</points>
<intersection>-21.5 2</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103,-20,103.5,-20</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>102,-21.5,103,-21.5</points>
<connection>
<GID>138</GID>
<name>OUT_5</name></connection>
<intersection>103 0</intersection></hsegment></shape></wire>
<wire>
<ID>984 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>241.5,-212,241.5,-212</points>
<connection>
<GID>620</GID>
<name>IN_0</name></connection>
<connection>
<GID>740</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>290 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-31,57,-30.5</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<connection>
<GID>49</GID>
<name>IN_B_1</name></connection></vsegment></shape></wire>
<wire>
<ID>654 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219,-126.5,219,-116.5</points>
<intersection>-126.5 2</intersection>
<intersection>-116.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>219,-116.5,220,-116.5</points>
<connection>
<GID>399</GID>
<name>IN_6</name></connection>
<intersection>219 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200.5,-126.5,219,-126.5</points>
<connection>
<GID>382</GID>
<name>OUT</name></connection>
<intersection>219 0</intersection></hsegment></shape></wire>
<wire>
<ID>291 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-32.5,57,-32</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<connection>
<GID>49</GID>
<name>IN_B_2</name></connection></vsegment></shape></wire>
<wire>
<ID>292 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-34.5,57,-33</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<connection>
<GID>49</GID>
<name>IN_B_3</name></connection></vsegment></shape></wire>
<wire>
<ID>289 </ID>
<shape>
<vsegment>
<ID>4</ID>
<points>65,-38,65,-36.5</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<connection>
<GID>49</GID>
<name>OUT_3</name></connection></vsegment></shape></wire>
<wire>
<ID>991 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>227,-115,227,-115</points>
<connection>
<GID>747</GID>
<name>IN_0</name></connection>
<connection>
<GID>399</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>616 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-113.5,142.5,-113.5</points>
<connection>
<GID>356</GID>
<name>IN_0</name></connection>
<connection>
<GID>368</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>983 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-206,245.5,-206</points>
<connection>
<GID>739</GID>
<name>IN_0</name></connection>
<connection>
<GID>605</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>936 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-166.5,138,-166.5</points>
<connection>
<GID>477</GID>
<name>IN_0</name></connection>
<connection>
<GID>691</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>876 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-58,194.5,-58</points>
<connection>
<GID>277</GID>
<name>IN_1</name></connection>
<connection>
<GID>629</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>715 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-166.5,142,-166.5</points>
<connection>
<GID>477</GID>
<name>OUT_0</name></connection>
<connection>
<GID>463</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>652 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>200.5,-114.5,220,-114.5</points>
<connection>
<GID>380</GID>
<name>OUT</name></connection>
<connection>
<GID>399</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>445 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-54,57,-54</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<connection>
<GID>79</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>447 </ID>
<shape>
<vsegment>
<ID>3</ID>
<points>57,-58,57,-56</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<connection>
<GID>71</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>753 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-138.5,245.5,-138.5</points>
<connection>
<GID>506</GID>
<name>IN_0</name></connection>
<connection>
<GID>514</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>448 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-60,57,-57</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<connection>
<GID>71</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>621 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-125.5,142.5,-125.5</points>
<connection>
<GID>359</GID>
<name>IN_0</name></connection>
<connection>
<GID>373</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>444 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-47,57,-45.5</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<connection>
<GID>71</GID>
<name>IN_B_0</name></connection></vsegment></shape></wire>
<wire>
<ID>441 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-48,57,-47.5</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<connection>
<GID>71</GID>
<name>IN_B_1</name></connection></vsegment></shape></wire>
<wire>
<ID>442 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-49.5,57,-49</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<connection>
<GID>71</GID>
<name>IN_B_2</name></connection></vsegment></shape></wire>
<wire>
<ID>443 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-51.5,57,-50</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<connection>
<GID>71</GID>
<name>IN_B_3</name></connection></vsegment></shape></wire>
<wire>
<ID>627 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167,-113.5,167,-108.5</points>
<intersection>-113.5 1</intersection>
<intersection>-108.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>167,-113.5,168,-113.5</points>
<connection>
<GID>376</GID>
<name>IN_2</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148.5,-108.5,167,-108.5</points>
<connection>
<GID>355</GID>
<name>OUT</name></connection>
<intersection>167 0</intersection></hsegment></shape></wire>
<wire>
<ID>478 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94,-32,94,-26.5</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-32,94,-32</points>
<connection>
<GID>134</GID>
<name>OUT_0</name></connection>
<intersection>94 0</intersection></hsegment></shape></wire>
<wire>
<ID>801 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-184,142,-184</points>
<connection>
<GID>557</GID>
<name>IN_0</name></connection>
<connection>
<GID>566</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>479 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93.5,-30,93.5,-25.5</points>
<intersection>-30 2</intersection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93.5,-25.5,94,-25.5</points>
<connection>
<GID>138</GID>
<name>IN_1</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-30,93.5,-30</points>
<connection>
<GID>134</GID>
<name>OUT_1</name></connection>
<intersection>93.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>810 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-210,142,-210</points>
<connection>
<GID>575</GID>
<name>IN_0</name></connection>
<connection>
<GID>563</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>657 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-93.5,246,-93.5</points>
<connection>
<GID>401</GID>
<name>IN_0</name></connection>
<connection>
<GID>409</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>480 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,-28,93,-24.5</points>
<intersection>-28 2</intersection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93,-24.5,94,-24.5</points>
<connection>
<GID>138</GID>
<name>IN_2</name></connection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-28,93,-28</points>
<connection>
<GID>134</GID>
<name>OUT_2</name></connection>
<intersection>93 0</intersection></hsegment></shape></wire>
<wire>
<ID>481 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92.5,-26,92.5,-23.5</points>
<intersection>-26 2</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92.5,-23.5,94,-23.5</points>
<connection>
<GID>138</GID>
<name>IN_3</name></connection>
<intersection>92.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-26,92.5,-26</points>
<connection>
<GID>134</GID>
<name>OUT_3</name></connection>
<intersection>92.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>485 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92.5,-22.5,92.5,-20</points>
<intersection>-22.5 1</intersection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92.5,-22.5,94,-22.5</points>
<connection>
<GID>138</GID>
<name>IN_4</name></connection>
<intersection>92.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-20,92.5,-20</points>
<connection>
<GID>130</GID>
<name>OUT_0</name></connection>
<intersection>92.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>484 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,-21.5,93,-18</points>
<intersection>-21.5 1</intersection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93,-21.5,94,-21.5</points>
<connection>
<GID>138</GID>
<name>IN_5</name></connection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-18,93,-18</points>
<connection>
<GID>130</GID>
<name>OUT_1</name></connection>
<intersection>93 0</intersection></hsegment></shape></wire>
<wire>
<ID>821 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167,-223,167,-208</points>
<intersection>-223 2</intersection>
<intersection>-208 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>148,-223,167,-223</points>
<connection>
<GID>565</GID>
<name>OUT</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>167,-208,167.5,-208</points>
<connection>
<GID>580</GID>
<name>IN_5</name></connection>
<intersection>167 0</intersection></hsegment></shape></wire>
<wire>
<ID>483 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93.5,-20.5,93.5,-16</points>
<intersection>-20.5 1</intersection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93.5,-20.5,94,-20.5</points>
<connection>
<GID>138</GID>
<name>IN_6</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-16,93.5,-16</points>
<connection>
<GID>130</GID>
<name>OUT_2</name></connection>
<intersection>93.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>519 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-64,142.5,-64</points>
<connection>
<GID>253</GID>
<name>IN_1</name></connection>
<connection>
<GID>264</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>482 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94,-19.5,94,-14</points>
<connection>
<GID>138</GID>
<name>IN_7</name></connection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-14,94,-14</points>
<connection>
<GID>130</GID>
<name>OUT_3</name></connection>
<intersection>94 0</intersection></hsegment></shape></wire>
<wire>
<ID>818 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167,-203,167,-193</points>
<intersection>-203 1</intersection>
<intersection>-193 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>167,-203,167.5,-203</points>
<connection>
<GID>580</GID>
<name>IN_1</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148,-193,167,-193</points>
<connection>
<GID>558</GID>
<name>OUT</name></connection>
<intersection>167 0</intersection></hsegment></shape></wire>
<wire>
<ID>488 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97,-28.5,97,-28.5</points>
<connection>
<GID>138</GID>
<name>clock</name></connection>
<connection>
<GID>158</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>489 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-30,102,-26.5</points>
<connection>
<GID>138</GID>
<name>OUT_0</name></connection>
<intersection>-30 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>102,-30,103.5,-30</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>102 0</intersection></hsegment></shape></wire>
<wire>
<ID>673 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271.5,-111.5,271.5,-95.5</points>
<connection>
<GID>424</GID>
<name>IN_0</name></connection>
<intersection>-95.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>252,-95.5,271.5,-95.5</points>
<connection>
<GID>401</GID>
<name>OUT</name></connection>
<intersection>271.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>496 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>102,-25.5,102.5,-25.5</points>
<connection>
<GID>138</GID>
<name>OUT_1</name></connection>
<intersection>102.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>102.5,-28,102.5,-25.5</points>
<intersection>-28 8</intersection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>102.5,-28,103.5,-28</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<intersection>102.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>817 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167.5,-202,167.5,-186</points>
<connection>
<GID>580</GID>
<name>IN_0</name></connection>
<intersection>-186 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>148,-186,167.5,-186</points>
<connection>
<GID>557</GID>
<name>OUT</name></connection>
<intersection>167.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>495 </ID>
<shape>
<vsegment>
<ID>5</ID>
<points>103,-26,103,-24.5</points>
<intersection>-26 8</intersection>
<intersection>-24.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>102,-24.5,103,-24.5</points>
<connection>
<GID>138</GID>
<name>OUT_2</name></connection>
<intersection>103 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>103,-26,103.5,-26</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<intersection>103 5</intersection></hsegment></shape></wire>
<wire>
<ID>515 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>142.5,-52,142.5,-52</points>
<connection>
<GID>251</GID>
<name>IN_2</name></connection>
<connection>
<GID>260</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>494 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>102,-24,103.5,-24</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<intersection>102 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>102,-24,102,-23.5</points>
<connection>
<GID>138</GID>
<name>OUT_3</name></connection>
<intersection>-24 5</intersection></vsegment></shape></wire>
<wire>
<ID>491 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-20.5,102.5,-18</points>
<intersection>-20.5 2</intersection>
<intersection>-18 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>102,-20.5,102.5,-20.5</points>
<connection>
<GID>138</GID>
<name>OUT_6</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>102.5,-18,103.5,-18</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>102.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>527 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-86,142.5,-86</points>
<connection>
<GID>272</GID>
<name>IN_0</name></connection>
<connection>
<GID>257</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>490 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-19.5,102,-16</points>
<connection>
<GID>138</GID>
<name>OUT_7</name></connection>
<intersection>-16 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>102,-16,103.5,-16</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>102 0</intersection></hsegment></shape></wire>
<wire>
<ID>710 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-152.5,142,-152.5</points>
<connection>
<GID>471</GID>
<name>IN_0</name></connection>
<connection>
<GID>460</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>719 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-176.5,142,-176.5</points>
<connection>
<GID>465</GID>
<name>IN_0</name></connection>
<connection>
<GID>462</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>938 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-178.5,142,-178.5</points>
<connection>
<GID>465</GID>
<name>IN_1</name></connection>
<connection>
<GID>693</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>878 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-70,194.5,-70</points>
<connection>
<GID>279</GID>
<name>IN_1</name></connection>
<connection>
<GID>631</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>725 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167,-177.5,167,-162.5</points>
<intersection>-177.5 2</intersection>
<intersection>-162.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>148,-177.5,167,-177.5</points>
<connection>
<GID>465</GID>
<name>OUT</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>167,-162.5,167.5,-162.5</points>
<connection>
<GID>481</GID>
<name>IN_5</name></connection>
<intersection>167 0</intersection></hsegment></shape></wire>
<wire>
<ID>734 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-152.5,194,-152.5</points>
<connection>
<GID>459</GID>
<name>IN_0</name></connection>
<connection>
<GID>493</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>942 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-154.5,194,-154.5</points>
<connection>
<GID>459</GID>
<name>IN_1</name></connection>
<connection>
<GID>698</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>780 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-192,90.5,-192</points>
<connection>
<GID>541</GID>
<name>IN_0</name></connection>
<connection>
<GID>532</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>747 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218.5,-158.5,218.5,-153.5</points>
<intersection>-158.5 1</intersection>
<intersection>-153.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218.5,-158.5,219.5,-158.5</points>
<connection>
<GID>504</GID>
<name>IN_2</name></connection>
<intersection>218.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200,-153.5,218.5,-153.5</points>
<connection>
<GID>459</GID>
<name>OUT</name></connection>
<intersection>218.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>501 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-66,116.5,-50</points>
<connection>
<GID>248</GID>
<name>IN_0</name></connection>
<intersection>-50 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>97,-50,116.5,-50</points>
<connection>
<GID>7</GID>
<name>OUT</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>708 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-146.5,142,-146.5</points>
<connection>
<GID>469</GID>
<name>IN_0</name></connection>
<connection>
<GID>458</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>505 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-119,116.5,-118.5</points>
<connection>
<GID>349</GID>
<name>IN_4</name></connection>
<connection>
<GID>231</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>712 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-158.5,142,-158.5</points>
<connection>
<GID>473</GID>
<name>IN_0</name></connection>
<connection>
<GID>461</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>874 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-50,194.5,-50</points>
<connection>
<GID>276</GID>
<name>IN_1</name></connection>
<connection>
<GID>627</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>721 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167.5,-156.5,167.5,-140.5</points>
<connection>
<GID>481</GID>
<name>IN_0</name></connection>
<intersection>-140.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>148,-140.5,167.5,-140.5</points>
<connection>
<GID>457</GID>
<name>OUT</name></connection>
<intersection>167.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>722 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167,-157.5,167,-147.5</points>
<intersection>-157.5 1</intersection>
<intersection>-147.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>167,-157.5,167.5,-157.5</points>
<connection>
<GID>481</GID>
<name>IN_1</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148,-147.5,167,-147.5</points>
<connection>
<GID>458</GID>
<name>OUT</name></connection>
<intersection>167 0</intersection></hsegment></shape></wire>
<wire>
<ID>884 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-52,246,-52</points>
<connection>
<GID>301</GID>
<name>IN_2</name></connection>
<connection>
<GID>637</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>723 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166.5,-158.5,166.5,-153.5</points>
<intersection>-158.5 1</intersection>
<intersection>-153.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166.5,-158.5,167.5,-158.5</points>
<connection>
<GID>481</GID>
<name>IN_2</name></connection>
<intersection>166.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148,-153.5,166.5,-153.5</points>
<connection>
<GID>460</GID>
<name>OUT</name></connection>
<intersection>166.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>724 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>148,-159.5,167.5,-159.5</points>
<connection>
<GID>461</GID>
<name>OUT</name></connection>
<connection>
<GID>481</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>331 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167.5,-164,167.5,-163.5</points>
<connection>
<GID>481</GID>
<name>IN_4</name></connection>
<connection>
<GID>222</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>726 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166.5,-171.5,166.5,-161.5</points>
<intersection>-171.5 2</intersection>
<intersection>-161.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166.5,-161.5,167.5,-161.5</points>
<connection>
<GID>481</GID>
<name>IN_6</name></connection>
<intersection>166.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148,-171.5,166.5,-171.5</points>
<connection>
<GID>464</GID>
<name>OUT</name></connection>
<intersection>166.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>727 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,-165.5,166,-160.5</points>
<intersection>-165.5 2</intersection>
<intersection>-160.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166,-160.5,167.5,-160.5</points>
<connection>
<GID>481</GID>
<name>IN_7</name></connection>
<intersection>166 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148,-165.5,166,-165.5</points>
<connection>
<GID>463</GID>
<name>OUT</name></connection>
<intersection>166 0</intersection></hsegment></shape></wire>
<wire>
<ID>994 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>174.5,-160,174.5,-160</points>
<connection>
<GID>481</GID>
<name>OUT</name></connection>
<connection>
<GID>750</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>736 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-158.5,194,-158.5</points>
<connection>
<GID>485</GID>
<name>IN_0</name></connection>
<connection>
<GID>495</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>943 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-160.5,194,-160.5</points>
<connection>
<GID>485</GID>
<name>IN_1</name></connection>
<connection>
<GID>699</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>748 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>200,-159.5,219.5,-159.5</points>
<connection>
<GID>485</GID>
<name>OUT</name></connection>
<connection>
<GID>504</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>612 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-101.5,142.5,-101.5</points>
<connection>
<GID>353</GID>
<name>IN_0</name></connection>
<connection>
<GID>364</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>963 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-186,142,-186</points>
<connection>
<GID>557</GID>
<name>IN_1</name></connection>
<connection>
<GID>719</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>964 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-188,142,-188</points>
<connection>
<GID>557</GID>
<name>IN_2</name></connection>
<connection>
<GID>720</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>640 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-113.5,194.5,-113.5</points>
<connection>
<GID>380</GID>
<name>IN_0</name></connection>
<connection>
<GID>390</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>544 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-68,194.5,-68</points>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<connection>
<GID>290</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>911 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-115.5,194.5,-115.5</points>
<connection>
<GID>380</GID>
<name>IN_1</name></connection>
<connection>
<GID>664</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>631 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166.5,-120.5,166.5,-115.5</points>
<intersection>-120.5 2</intersection>
<intersection>-115.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166.5,-115.5,168,-115.5</points>
<connection>
<GID>376</GID>
<name>IN_7</name></connection>
<intersection>166.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148.5,-120.5,166.5,-120.5</points>
<connection>
<GID>358</GID>
<name>OUT</name></connection>
<intersection>166.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>466 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-48,91,-48</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<connection>
<GID>142</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>467 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-50,91,-50</points>
<connection>
<GID>7</GID>
<name>IN_1</name></connection>
<connection>
<GID>146</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>798 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-217,115,-207</points>
<intersection>-217 2</intersection>
<intersection>-207 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,-207,116,-207</points>
<connection>
<GID>554</GID>
<name>IN_6</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>96.5,-217,115,-217</points>
<connection>
<GID>536</GID>
<name>OUT</name></connection>
<intersection>115 0</intersection></hsegment></shape></wire>
<wire>
<ID>645 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-125.5,194.5,-125.5</points>
<connection>
<GID>382</GID>
<name>IN_0</name></connection>
<connection>
<GID>395</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>468 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>91,-52,91,-52</points>
<connection>
<GID>7</GID>
<name>IN_2</name></connection>
<connection>
<GID>150</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>469 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-56,91,-56</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<connection>
<GID>154</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>619 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-121.5,142.5,-121.5</points>
<connection>
<GID>358</GID>
<name>IN_1</name></connection>
<connection>
<GID>372</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>470 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-58,91,-58</points>
<connection>
<GID>36</GID>
<name>IN_1</name></connection>
<connection>
<GID>160</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>523 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-76,142.5,-76</points>
<connection>
<GID>255</GID>
<name>IN_1</name></connection>
<connection>
<GID>269</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>502 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116,-67,116,-57</points>
<intersection>-67 1</intersection>
<intersection>-57 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116,-67,116.5,-67</points>
<connection>
<GID>248</GID>
<name>IN_1</name></connection>
<intersection>116 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97,-57,116,-57</points>
<connection>
<GID>36</GID>
<name>OUT</name></connection>
<intersection>116 0</intersection></hsegment></shape></wire>
<wire>
<ID>894 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-109.5,91,-109.5</points>
<connection>
<GID>328</GID>
<name>IN_1</name></connection>
<connection>
<GID>647</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>741 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-170.5,194,-170.5</points>
<connection>
<GID>487</GID>
<name>IN_0</name></connection>
<connection>
<GID>500</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>945 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-172.5,194,-172.5</points>
<connection>
<GID>487</GID>
<name>IN_1</name></connection>
<connection>
<GID>701</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>750 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218.5,-171.5,218.5,-161.5</points>
<intersection>-171.5 2</intersection>
<intersection>-161.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218.5,-161.5,219.5,-161.5</points>
<connection>
<GID>504</GID>
<name>IN_6</name></connection>
<intersection>218.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200,-171.5,218.5,-171.5</points>
<connection>
<GID>487</GID>
<name>OUT</name></connection>
<intersection>218.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>473 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-62,91,-62</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<connection>
<GID>226</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>474 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-64,91,-64</points>
<connection>
<GID>120</GID>
<name>IN_1</name></connection>
<connection>
<GID>228</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>825 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-184,194,-184</points>
<connection>
<GID>582</GID>
<name>IN_0</name></connection>
<connection>
<GID>587</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>503 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-68,115.5,-63</points>
<intersection>-68 1</intersection>
<intersection>-63 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115.5,-68,116.5,-68</points>
<connection>
<GID>248</GID>
<name>IN_2</name></connection>
<intersection>115.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97,-63,115.5,-63</points>
<connection>
<GID>120</GID>
<name>OUT</name></connection>
<intersection>115.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>714 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-164.5,142,-164.5</points>
<connection>
<GID>475</GID>
<name>IN_0</name></connection>
<connection>
<GID>463</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>813 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-216,142,-216</points>
<connection>
<GID>564</GID>
<name>IN_0</name></connection>
<connection>
<GID>578</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>475 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-68,91,-68</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<connection>
<GID>230</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>806 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-198,142,-198</points>
<connection>
<GID>571</GID>
<name>IN_0</name></connection>
<connection>
<GID>560</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>653 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219.5,-132.5,219.5,-117.5</points>
<intersection>-132.5 2</intersection>
<intersection>-117.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>200.5,-132.5,219.5,-132.5</points>
<connection>
<GID>383</GID>
<name>OUT</name></connection>
<intersection>219.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>219.5,-117.5,220,-117.5</points>
<connection>
<GID>399</GID>
<name>IN_5</name></connection>
<intersection>219.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>476 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-70,91,-70</points>
<connection>
<GID>124</GID>
<name>IN_1</name></connection>
<connection>
<GID>232</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>508 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>97,-69,116.5,-69</points>
<connection>
<GID>124</GID>
<name>OUT</name></connection>
<connection>
<GID>248</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>477 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-74,91,-74</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<connection>
<GID>234</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>487 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-76,91,-76</points>
<connection>
<GID>128</GID>
<name>IN_1</name></connection>
<connection>
<GID>238</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>511 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-75,115,-70</points>
<intersection>-75 2</intersection>
<intersection>-70 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,-70,116.5,-70</points>
<connection>
<GID>248</GID>
<name>IN_7</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97,-75,115,-75</points>
<connection>
<GID>128</GID>
<name>OUT</name></connection>
<intersection>115 0</intersection></hsegment></shape></wire>
<wire>
<ID>493 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-80,91,-80</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<connection>
<GID>240</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>535 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166.5,-75,166.5,-70</points>
<intersection>-75 2</intersection>
<intersection>-70 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166.5,-70,168,-70</points>
<connection>
<GID>274</GID>
<name>IN_7</name></connection>
<intersection>166.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148.5,-75,166.5,-75</points>
<connection>
<GID>255</GID>
<name>OUT</name></connection>
<intersection>166.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>498 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-82,91,-82</points>
<connection>
<GID>132</GID>
<name>IN_1</name></connection>
<connection>
<GID>242</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>531 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167,-68,167,-63</points>
<intersection>-68 1</intersection>
<intersection>-63 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>167,-68,168,-68</points>
<connection>
<GID>274</GID>
<name>IN_2</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148.5,-63,167,-63</points>
<connection>
<GID>253</GID>
<name>OUT</name></connection>
<intersection>167 0</intersection></hsegment></shape></wire>
<wire>
<ID>510 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-81,115.5,-71</points>
<intersection>-81 2</intersection>
<intersection>-71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115.5,-71,116.5,-71</points>
<connection>
<GID>248</GID>
<name>IN_6</name></connection>
<intersection>115.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97,-81,115.5,-81</points>
<connection>
<GID>132</GID>
<name>OUT</name></connection>
<intersection>115.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>499 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-86,91,-86</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<connection>
<GID>244</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>525 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-80,142.5,-80</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<connection>
<GID>270</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>348 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>90,-88,91,-88</points>
<connection>
<GID>243</GID>
<name>OUT_0</name></connection>
<connection>
<GID>136</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>509 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116,-87,116,-72</points>
<intersection>-87 2</intersection>
<intersection>-72 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>97,-87,116,-87</points>
<connection>
<GID>136</GID>
<name>OUT</name></connection>
<intersection>116 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>116,-72,116.5,-72</points>
<connection>
<GID>248</GID>
<name>IN_5</name></connection>
<intersection>116 0</intersection></hsegment></shape></wire>
<wire>
<ID>643 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-121.5,194.5,-121.5</points>
<connection>
<GID>381</GID>
<name>IN_1</name></connection>
<connection>
<GID>394</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>804 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-192,142,-192</points>
<connection>
<GID>558</GID>
<name>IN_0</name></connection>
<connection>
<GID>569</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>606 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-126.5,115.5,-116.5</points>
<intersection>-126.5 2</intersection>
<intersection>-116.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115.5,-116.5,116.5,-116.5</points>
<connection>
<GID>349</GID>
<name>IN_6</name></connection>
<intersection>115.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97,-126.5,115.5,-126.5</points>
<connection>
<GID>331</GID>
<name>OUT</name></connection>
<intersection>115.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>965 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-194,142,-194</points>
<connection>
<GID>558</GID>
<name>IN_1</name></connection>
<connection>
<GID>721</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>815 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-222,142,-222</points>
<connection>
<GID>562</GID>
<name>IN_0</name></connection>
<connection>
<GID>565</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>669 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-125.5,246,-125.5</points>
<connection>
<GID>407</GID>
<name>IN_0</name></connection>
<connection>
<GID>421</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>822 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166.5,-217,166.5,-207</points>
<intersection>-217 2</intersection>
<intersection>-207 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166.5,-207,167.5,-207</points>
<connection>
<GID>580</GID>
<name>IN_6</name></connection>
<intersection>166.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148,-217,166.5,-217</points>
<connection>
<GID>564</GID>
<name>OUT</name></connection>
<intersection>166.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>492 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-76,87,-76</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<connection>
<GID>238</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>903 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-115.5,142.5,-115.5</points>
<connection>
<GID>656</GID>
<name>IN_0</name></connection>
<connection>
<GID>356</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>536 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-73.5,116.5,-73</points>
<connection>
<GID>248</GID>
<name>IN_4</name></connection>
<connection>
<GID>239</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>512 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>123.5,-69.5,123.5,-69.5</points>
<connection>
<GID>248</GID>
<name>OUT</name></connection>
<connection>
<GID>250</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>513 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-48,142.5,-48</points>
<connection>
<GID>251</GID>
<name>IN_0</name></connection>
<connection>
<GID>258</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>514 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-50,142.5,-50</points>
<connection>
<GID>251</GID>
<name>IN_1</name></connection>
<connection>
<GID>259</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>529 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168,-66,168,-50</points>
<connection>
<GID>274</GID>
<name>IN_0</name></connection>
<intersection>-50 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>148.5,-50,168,-50</points>
<connection>
<GID>251</GID>
<name>OUT</name></connection>
<intersection>168 0</intersection></hsegment></shape></wire>
<wire>
<ID>517 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>142.5,-58,142.5,-58</points>
<connection>
<GID>252</GID>
<name>IN_1</name></connection>
<connection>
<GID>262</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>530 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167.5,-67,167.5,-57</points>
<intersection>-67 1</intersection>
<intersection>-57 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>167.5,-67,168,-67</points>
<connection>
<GID>274</GID>
<name>IN_1</name></connection>
<intersection>167.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148.5,-57,167.5,-57</points>
<connection>
<GID>252</GID>
<name>OUT</name></connection>
<intersection>167.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>901 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-103.5,142.5,-103.5</points>
<connection>
<GID>353</GID>
<name>IN_1</name></connection>
<connection>
<GID>654</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>542 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-62,194.5,-62</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<connection>
<GID>288</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>877 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-64,194.5,-64</points>
<connection>
<GID>278</GID>
<name>IN_1</name></connection>
<connection>
<GID>630</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>555 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219,-68,219,-63</points>
<intersection>-68 1</intersection>
<intersection>-63 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>219,-68,220,-68</points>
<connection>
<GID>299</GID>
<name>IN_2</name></connection>
<intersection>219 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200.5,-63,219,-63</points>
<connection>
<GID>278</GID>
<name>OUT</name></connection>
<intersection>219 0</intersection></hsegment></shape></wire>
<wire>
<ID>518 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-62,142.5,-62</points>
<connection>
<GID>253</GID>
<name>IN_0</name></connection>
<connection>
<GID>263</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>520 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-68,142.5,-68</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<connection>
<GID>265</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>521 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-70,142.5,-70</points>
<connection>
<GID>254</GID>
<name>IN_1</name></connection>
<connection>
<GID>266</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>532 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>148.5,-69,168,-69</points>
<connection>
<GID>274</GID>
<name>IN_3</name></connection>
<connection>
<GID>254</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>522 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-74,142.5,-74</points>
<connection>
<GID>255</GID>
<name>IN_0</name></connection>
<connection>
<GID>267</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>808 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-204,142,-204</points>
<connection>
<GID>561</GID>
<name>IN_0</name></connection>
<connection>
<GID>573</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>820 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>148,-205,167.5,-205</points>
<connection>
<GID>561</GID>
<name>OUT</name></connection>
<connection>
<GID>580</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>526 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-82,142.5,-82</points>
<connection>
<GID>256</GID>
<name>IN_1</name></connection>
<connection>
<GID>271</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>534 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167,-81,167,-71</points>
<intersection>-81 2</intersection>
<intersection>-71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>167,-71,168,-71</points>
<connection>
<GID>274</GID>
<name>IN_6</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148.5,-81,167,-81</points>
<connection>
<GID>256</GID>
<name>OUT</name></connection>
<intersection>167 0</intersection></hsegment></shape></wire>
<wire>
<ID>832 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-204,194,-204</points>
<connection>
<GID>592</GID>
<name>IN_0</name></connection>
<connection>
<GID>428</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>881 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-88,142.5,-88</points>
<connection>
<GID>257</GID>
<name>IN_1</name></connection>
<connection>
<GID>634</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>533 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167.5,-87,167.5,-72</points>
<intersection>-87 2</intersection>
<intersection>-72 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>148.5,-87,167.5,-87</points>
<connection>
<GID>257</GID>
<name>OUT</name></connection>
<intersection>167.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>167.5,-72,168,-72</points>
<connection>
<GID>274</GID>
<name>IN_5</name></connection>
<intersection>167.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>506 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271.5,-73.5,271.5,-73</points>
<connection>
<GID>324</GID>
<name>IN_4</name></connection>
<connection>
<GID>233</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>677 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271,-132.5,271,-117.5</points>
<intersection>-132.5 2</intersection>
<intersection>-117.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>252,-132.5,271,-132.5</points>
<connection>
<GID>408</GID>
<name>OUT</name></connection>
<intersection>271 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>271,-117.5,271.5,-117.5</points>
<connection>
<GID>424</GID>
<name>IN_5</name></connection>
<intersection>271 0</intersection></hsegment></shape></wire>
<wire>
<ID>830 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-198,194,-198</points>
<connection>
<GID>559</GID>
<name>IN_0</name></connection>
<connection>
<GID>590</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>500 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>220,-119,220,-118.5</points>
<connection>
<GID>399</GID>
<name>IN_4</name></connection>
<connection>
<GID>227</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>970 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-224,142,-224</points>
<connection>
<GID>565</GID>
<name>IN_1</name></connection>
<connection>
<GID>726</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>837 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-216,194,-216</points>
<connection>
<GID>596</GID>
<name>IN_0</name></connection>
<connection>
<GID>585</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>528 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168,-73.5,168,-73</points>
<connection>
<GID>274</GID>
<name>IN_4</name></connection>
<connection>
<GID>237</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>982 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-200,245.5,-200</points>
<connection>
<GID>738</GID>
<name>IN_0</name></connection>
<connection>
<GID>604</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>841 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219.5,-202,219.5,-186</points>
<connection>
<GID>600</GID>
<name>IN_0</name></connection>
<intersection>-186 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>200,-186,219.5,-186</points>
<connection>
<GID>582</GID>
<name>OUT</name></connection>
<intersection>219.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>842 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219,-203,219,-193</points>
<intersection>-203 1</intersection>
<intersection>-193 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>219,-203,219.5,-203</points>
<connection>
<GID>600</GID>
<name>IN_1</name></connection>
<intersection>219 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200,-193,219,-193</points>
<connection>
<GID>583</GID>
<name>OUT</name></connection>
<intersection>219 0</intersection></hsegment></shape></wire>
<wire>
<ID>843 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218.5,-204,218.5,-199</points>
<intersection>-204 1</intersection>
<intersection>-199 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218.5,-204,219.5,-204</points>
<connection>
<GID>600</GID>
<name>IN_2</name></connection>
<intersection>218.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200,-199,218.5,-199</points>
<connection>
<GID>559</GID>
<name>OUT</name></connection>
<intersection>218.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>844 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>200,-205,219.5,-205</points>
<connection>
<GID>428</GID>
<name>OUT</name></connection>
<connection>
<GID>600</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>793 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116,-202,116,-186</points>
<connection>
<GID>554</GID>
<name>IN_0</name></connection>
<intersection>-186 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>96.5,-186,116,-186</points>
<connection>
<GID>531</GID>
<name>OUT</name></connection>
<intersection>116 0</intersection></hsegment></shape></wire>
<wire>
<ID>471 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219.5,-164,219.5,-163.5</points>
<connection>
<GID>504</GID>
<name>IN_4</name></connection>
<connection>
<GID>223</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>104 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219.5,-209.5,219.5,-209</points>
<connection>
<GID>600</GID>
<name>IN_4</name></connection>
<connection>
<GID>148</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>845 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219,-223,219,-208</points>
<intersection>-223 2</intersection>
<intersection>-208 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>200,-223,219,-223</points>
<connection>
<GID>586</GID>
<name>OUT</name></connection>
<intersection>219 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>219,-208,219.5,-208</points>
<connection>
<GID>600</GID>
<name>IN_5</name></connection>
<intersection>219 0</intersection></hsegment></shape></wire>
<wire>
<ID>846 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218.5,-217,218.5,-207</points>
<intersection>-217 2</intersection>
<intersection>-207 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218.5,-207,219.5,-207</points>
<connection>
<GID>600</GID>
<name>IN_6</name></connection>
<intersection>218.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200,-217,218.5,-217</points>
<connection>
<GID>585</GID>
<name>OUT</name></connection>
<intersection>218.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>847 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218,-211,218,-206</points>
<intersection>-211 2</intersection>
<intersection>-206 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218,-206,219.5,-206</points>
<connection>
<GID>600</GID>
<name>IN_7</name></connection>
<intersection>218 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200,-211,218,-211</points>
<connection>
<GID>584</GID>
<name>OUT</name></connection>
<intersection>218 0</intersection></hsegment></shape></wire>
<wire>
<ID>507 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>220,-73.5,220,-73</points>
<connection>
<GID>299</GID>
<name>IN_4</name></connection>
<connection>
<GID>235</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>524 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,-76,138.5,-76</points>
<connection>
<GID>268</GID>
<name>IN_0</name></connection>
<connection>
<GID>269</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>854 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-198,245.5,-198</points>
<connection>
<GID>604</GID>
<name>IN_0</name></connection>
<connection>
<GID>614</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>867 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270,-204,270,-199</points>
<intersection>-204 1</intersection>
<intersection>-199 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>270,-204,271,-204</points>
<connection>
<GID>624</GID>
<name>IN_2</name></connection>
<intersection>270 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>251.5,-199,270,-199</points>
<connection>
<GID>604</GID>
<name>OUT</name></connection>
<intersection>270 0</intersection></hsegment></shape></wire>
<wire>
<ID>990 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>175,-115,175,-115</points>
<connection>
<GID>746</GID>
<name>IN_0</name></connection>
<connection>
<GID>376</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>861 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-216,245.5,-216</points>
<connection>
<GID>608</GID>
<name>IN_0</name></connection>
<connection>
<GID>621</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>862 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-218,245.5,-218</points>
<connection>
<GID>608</GID>
<name>IN_1</name></connection>
<connection>
<GID>622</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>717 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-170.5,142,-170.5</points>
<connection>
<GID>464</GID>
<name>IN_0</name></connection>
<connection>
<GID>478</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>870 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270,-217,270,-207</points>
<intersection>-217 2</intersection>
<intersection>-207 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>270,-207,271,-207</points>
<connection>
<GID>624</GID>
<name>IN_6</name></connection>
<intersection>270 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>251.5,-217,270,-217</points>
<connection>
<GID>608</GID>
<name>OUT</name></connection>
<intersection>270 0</intersection></hsegment></shape></wire>
<wire>
<ID>986 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>175,-69.5,175,-69.5</points>
<connection>
<GID>274</GID>
<name>OUT</name></connection>
<connection>
<GID>742</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>537 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-48,194.5,-48</points>
<connection>
<GID>276</GID>
<name>IN_0</name></connection>
<connection>
<GID>283</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>875 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-52,194.5,-52</points>
<connection>
<GID>276</GID>
<name>IN_2</name></connection>
<connection>
<GID>628</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>553 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>220,-66,220,-50</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<intersection>-50 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>200.5,-50,220,-50</points>
<connection>
<GID>276</GID>
<name>OUT</name></connection>
<intersection>220 0</intersection></hsegment></shape></wire>
<wire>
<ID>540 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-56,194.5,-56</points>
<connection>
<GID>277</GID>
<name>IN_0</name></connection>
<connection>
<GID>286</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>913 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-127.5,194.5,-127.5</points>
<connection>
<GID>382</GID>
<name>IN_1</name></connection>
<connection>
<GID>666</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>554 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219.5,-67,219.5,-57</points>
<intersection>-67 1</intersection>
<intersection>-57 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>219.5,-67,220,-67</points>
<connection>
<GID>299</GID>
<name>IN_1</name></connection>
<intersection>219.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200.5,-57,219.5,-57</points>
<connection>
<GID>277</GID>
<name>OUT</name></connection>
<intersection>219.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>998 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>174.5,-205.5,174.5,-205.5</points>
<connection>
<GID>754</GID>
<name>IN_0</name></connection>
<connection>
<GID>580</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>907 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-95.5,194.5,-95.5</points>
<connection>
<GID>660</GID>
<name>IN_0</name></connection>
<connection>
<GID>378</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>556 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>200.5,-69,220,-69</points>
<connection>
<GID>279</GID>
<name>OUT</name></connection>
<connection>
<GID>299</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>905 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-127.5,142.5,-127.5</points>
<connection>
<GID>359</GID>
<name>IN_1</name></connection>
<connection>
<GID>658</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>546 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-74,194.5,-74</points>
<connection>
<GID>280</GID>
<name>IN_0</name></connection>
<connection>
<GID>292</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>547 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-76,194.5,-76</points>
<connection>
<GID>280</GID>
<name>IN_1</name></connection>
<connection>
<GID>294</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>559 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218.5,-75,218.5,-70</points>
<intersection>-75 2</intersection>
<intersection>-70 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218.5,-70,220,-70</points>
<connection>
<GID>299</GID>
<name>IN_7</name></connection>
<intersection>218.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200.5,-75,218.5,-75</points>
<connection>
<GID>280</GID>
<name>OUT</name></connection>
<intersection>218.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>856 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-204,245.5,-204</points>
<connection>
<GID>616</GID>
<name>IN_0</name></connection>
<connection>
<GID>605</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>549 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-80,194.5,-80</points>
<connection>
<GID>281</GID>
<name>IN_0</name></connection>
<connection>
<GID>295</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>880 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-82,194.5,-82</points>
<connection>
<GID>281</GID>
<name>IN_1</name></connection>
<connection>
<GID>633</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>917 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-103.5,246,-103.5</points>
<connection>
<GID>670</GID>
<name>IN_0</name></connection>
<connection>
<GID>402</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>558 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219,-81,219,-71</points>
<intersection>-81 2</intersection>
<intersection>-71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>219,-71,220,-71</points>
<connection>
<GID>299</GID>
<name>IN_6</name></connection>
<intersection>219 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200.5,-81,219,-81</points>
<connection>
<GID>281</GID>
<name>OUT</name></connection>
<intersection>219 0</intersection></hsegment></shape></wire>
<wire>
<ID>551 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-86,194.5,-86</points>
<connection>
<GID>282</GID>
<name>IN_0</name></connection>
<connection>
<GID>297</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>729 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-138.5,194,-138.5</points>
<connection>
<GID>483</GID>
<name>IN_0</name></connection>
<connection>
<GID>489</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>882 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-88,194.5,-88</points>
<connection>
<GID>282</GID>
<name>IN_1</name></connection>
<connection>
<GID>635</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>557 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219.5,-87,219.5,-72</points>
<intersection>-87 2</intersection>
<intersection>-72 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>200.5,-87,219.5,-87</points>
<connection>
<GID>282</GID>
<name>OUT</name></connection>
<intersection>219.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>219.5,-72,220,-72</points>
<connection>
<GID>299</GID>
<name>IN_5</name></connection>
<intersection>219.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>859 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-212,245.5,-212</points>
<connection>
<GID>620</GID>
<name>OUT_0</name></connection>
<connection>
<GID>607</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>865 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271,-202,271,-186</points>
<connection>
<GID>624</GID>
<name>IN_0</name></connection>
<intersection>-186 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>251.5,-186,271,-186</points>
<connection>
<GID>602</GID>
<name>OUT</name></connection>
<intersection>271 0</intersection></hsegment></shape></wire>
<wire>
<ID>866 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,-203,270.5,-193</points>
<intersection>-203 1</intersection>
<intersection>-193 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>270.5,-203,271,-203</points>
<connection>
<GID>624</GID>
<name>IN_1</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>251.5,-193,270.5,-193</points>
<connection>
<GID>603</GID>
<name>OUT</name></connection>
<intersection>270.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>868 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>251.5,-205,271,-205</points>
<connection>
<GID>605</GID>
<name>OUT</name></connection>
<connection>
<GID>624</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>869 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,-223,270.5,-208</points>
<intersection>-223 2</intersection>
<intersection>-208 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>251.5,-223,270.5,-223</points>
<connection>
<GID>609</GID>
<name>OUT</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>270.5,-208,271,-208</points>
<connection>
<GID>624</GID>
<name>IN_5</name></connection>
<intersection>270.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>871 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269.5,-211,269.5,-206</points>
<intersection>-211 2</intersection>
<intersection>-206 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>269.5,-206,271,-206</points>
<connection>
<GID>624</GID>
<name>IN_7</name></connection>
<intersection>269.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>251.5,-211,269.5,-211</points>
<connection>
<GID>607</GID>
<name>OUT</name></connection>
<intersection>269.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1000 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278,-205.5,278,-205.5</points>
<connection>
<GID>624</GID>
<name>OUT</name></connection>
<connection>
<GID>756</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>879 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190.5,-76,190.5,-76</points>
<connection>
<GID>294</GID>
<name>IN_0</name></connection>
<connection>
<GID>632</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>909 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-103.5,194.5,-103.5</points>
<connection>
<GID>662</GID>
<name>IN_0</name></connection>
<connection>
<GID>379</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>883 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-50,246,-50</points>
<connection>
<GID>636</GID>
<name>IN_0</name></connection>
<connection>
<GID>301</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>561 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-48,246,-48</points>
<connection>
<GID>301</GID>
<name>IN_0</name></connection>
<connection>
<GID>309</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>577 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271.5,-66,271.5,-50</points>
<connection>
<GID>324</GID>
<name>IN_0</name></connection>
<intersection>-50 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>252,-50,271.5,-50</points>
<connection>
<GID>301</GID>
<name>OUT</name></connection>
<intersection>271.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>915 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-95.5,246,-95.5</points>
<connection>
<GID>668</GID>
<name>IN_0</name></connection>
<connection>
<GID>401</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>564 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-56,246,-56</points>
<connection>
<GID>302</GID>
<name>IN_0</name></connection>
<connection>
<GID>312</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>885 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-58,246,-58</points>
<connection>
<GID>302</GID>
<name>IN_1</name></connection>
<connection>
<GID>638</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>578 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271,-67,271,-57</points>
<intersection>-67 1</intersection>
<intersection>-57 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>271,-67,271.5,-67</points>
<connection>
<GID>324</GID>
<name>IN_1</name></connection>
<intersection>271 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>252,-57,271,-57</points>
<connection>
<GID>302</GID>
<name>OUT</name></connection>
<intersection>271 0</intersection></hsegment></shape></wire>
<wire>
<ID>897 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-127.5,91,-127.5</points>
<connection>
<GID>650</GID>
<name>IN_0</name></connection>
<connection>
<GID>331</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>925 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-148.5,90.5,-148.5</points>
<connection>
<GID>432</GID>
<name>IN_1</name></connection>
<connection>
<GID>678</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>566 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-62,246,-62</points>
<connection>
<GID>303</GID>
<name>IN_0</name></connection>
<connection>
<GID>314</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>886 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-64,246,-64</points>
<connection>
<GID>303</GID>
<name>IN_1</name></connection>
<connection>
<GID>639</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>579 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,-68,270.5,-63</points>
<intersection>-68 1</intersection>
<intersection>-63 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>270.5,-68,271.5,-68</points>
<connection>
<GID>324</GID>
<name>IN_2</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>252,-63,270.5,-63</points>
<connection>
<GID>303</GID>
<name>OUT</name></connection>
<intersection>270.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>935 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-160.5,142,-160.5</points>
<connection>
<GID>461</GID>
<name>IN_1</name></connection>
<connection>
<GID>690</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>568 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-68,246,-68</points>
<connection>
<GID>304</GID>
<name>IN_0</name></connection>
<connection>
<GID>316</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>887 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-70,246,-70</points>
<connection>
<GID>304</GID>
<name>IN_1</name></connection>
<connection>
<GID>640</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>580 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>252,-69,271.5,-69</points>
<connection>
<GID>304</GID>
<name>OUT</name></connection>
<connection>
<GID>324</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>953 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-172.5,245.5,-172.5</points>
<connection>
<GID>512</GID>
<name>IN_1</name></connection>
<connection>
<GID>709</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>749 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219,-177.5,219,-162.5</points>
<intersection>-177.5 2</intersection>
<intersection>-162.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>200,-177.5,219,-177.5</points>
<connection>
<GID>488</GID>
<name>OUT</name></connection>
<intersection>219 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>219,-162.5,219.5,-162.5</points>
<connection>
<GID>504</GID>
<name>IN_5</name></connection>
<intersection>219 0</intersection></hsegment></shape></wire>
<wire>
<ID>774 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270,-171.5,270,-161.5</points>
<intersection>-171.5 2</intersection>
<intersection>-161.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>270,-161.5,271,-161.5</points>
<connection>
<GID>529</GID>
<name>IN_6</name></connection>
<intersection>270 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>251.5,-171.5,270,-171.5</points>
<connection>
<GID>512</GID>
<name>OUT</name></connection>
<intersection>270 0</intersection></hsegment></shape></wire>
<wire>
<ID>575 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-86,246,-86</points>
<connection>
<GID>305</GID>
<name>IN_0</name></connection>
<connection>
<GID>308</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>929 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-172.5,90.5,-172.5</points>
<connection>
<GID>436</GID>
<name>IN_1</name></connection>
<connection>
<GID>682</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>570 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-74,246,-74</points>
<connection>
<GID>306</GID>
<name>IN_0</name></connection>
<connection>
<GID>318</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>571 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-76,246,-76</points>
<connection>
<GID>306</GID>
<name>IN_1</name></connection>
<connection>
<GID>320</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>583 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270,-75,270,-70</points>
<intersection>-75 2</intersection>
<intersection>-70 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>270,-70,271.5,-70</points>
<connection>
<GID>324</GID>
<name>IN_7</name></connection>
<intersection>270 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>252,-75,270,-75</points>
<connection>
<GID>306</GID>
<name>OUT</name></connection>
<intersection>270 0</intersection></hsegment></shape></wire>
<wire>
<ID>573 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-80,246,-80</points>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<connection>
<GID>321</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>582 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,-81,270.5,-71</points>
<intersection>-81 2</intersection>
<intersection>-71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>270.5,-71,271.5,-71</points>
<connection>
<GID>324</GID>
<name>IN_6</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>252,-81,270.5,-81</points>
<connection>
<GID>307</GID>
<name>OUT</name></connection>
<intersection>270.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>890 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-88,246,-88</points>
<connection>
<GID>308</GID>
<name>IN_1</name></connection>
<connection>
<GID>643</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>581 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271,-87,271,-72</points>
<intersection>-87 2</intersection>
<intersection>-72 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>252,-87,271,-87</points>
<connection>
<GID>308</GID>
<name>OUT</name></connection>
<intersection>271 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>271,-72,271.5,-72</points>
<connection>
<GID>324</GID>
<name>IN_5</name></connection>
<intersection>271 0</intersection></hsegment></shape></wire>
<wire>
<ID>743 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-176.5,194,-176.5</points>
<connection>
<GID>488</GID>
<name>IN_0</name></connection>
<connection>
<GID>502</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>888 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242,-76,242,-76</points>
<connection>
<GID>320</GID>
<name>IN_0</name></connection>
<connection>
<GID>641</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>585 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-93.5,91,-93.5</points>
<connection>
<GID>326</GID>
<name>IN_0</name></connection>
<connection>
<GID>333</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>891 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-95.5,91,-95.5</points>
<connection>
<GID>326</GID>
<name>IN_1</name></connection>
<connection>
<GID>644</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>892 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-97.5,91,-97.5</points>
<connection>
<GID>326</GID>
<name>IN_2</name></connection>
<connection>
<GID>645</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>601 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-111.5,116.5,-95.5</points>
<connection>
<GID>349</GID>
<name>IN_0</name></connection>
<intersection>-95.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>97,-95.5,116.5,-95.5</points>
<connection>
<GID>326</GID>
<name>OUT</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>588 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-101.5,91,-101.5</points>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<connection>
<GID>336</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>961 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-218,90.5,-218</points>
<connection>
<GID>536</GID>
<name>IN_1</name></connection>
<connection>
<GID>717</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>602 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116,-112.5,116,-102.5</points>
<intersection>-112.5 1</intersection>
<intersection>-102.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116,-112.5,116.5,-112.5</points>
<connection>
<GID>349</GID>
<name>IN_1</name></connection>
<intersection>116 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97,-102.5,116,-102.5</points>
<connection>
<GID>327</GID>
<name>OUT</name></connection>
<intersection>116 0</intersection></hsegment></shape></wire>
<wire>
<ID>590 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-107.5,91,-107.5</points>
<connection>
<GID>328</GID>
<name>IN_0</name></connection>
<connection>
<GID>338</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>592 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-113.5,91,-113.5</points>
<connection>
<GID>329</GID>
<name>IN_0</name></connection>
<connection>
<GID>340</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>895 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-115.5,91,-115.5</points>
<connection>
<GID>329</GID>
<name>IN_1</name></connection>
<connection>
<GID>648</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>604 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>97,-114.5,116.5,-114.5</points>
<connection>
<GID>329</GID>
<name>OUT</name></connection>
<connection>
<GID>349</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>594 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-119.5,91,-119.5</points>
<connection>
<GID>330</GID>
<name>IN_0</name></connection>
<connection>
<GID>342</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>595 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-121.5,91,-121.5</points>
<connection>
<GID>330</GID>
<name>IN_1</name></connection>
<connection>
<GID>344</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>607 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-120.5,115,-115.5</points>
<intersection>-120.5 2</intersection>
<intersection>-115.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,-115.5,116.5,-115.5</points>
<connection>
<GID>349</GID>
<name>IN_7</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97,-120.5,115,-120.5</points>
<connection>
<GID>330</GID>
<name>OUT</name></connection>
<intersection>115 0</intersection></hsegment></shape></wire>
<wire>
<ID>597 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>91,-125.5,91,-125.5</points>
<connection>
<GID>331</GID>
<name>IN_0</name></connection>
<connection>
<GID>345</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>599 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-131.5,91,-131.5</points>
<connection>
<GID>332</GID>
<name>IN_0</name></connection>
<connection>
<GID>347</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>898 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-133.5,91,-133.5</points>
<connection>
<GID>332</GID>
<name>IN_1</name></connection>
<connection>
<GID>651</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>605 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116,-132.5,116,-117.5</points>
<intersection>-132.5 2</intersection>
<intersection>-117.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>97,-132.5,116,-132.5</points>
<connection>
<GID>332</GID>
<name>OUT</name></connection>
<intersection>116 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>116,-117.5,116.5,-117.5</points>
<connection>
<GID>349</GID>
<name>IN_5</name></connection>
<intersection>116 0</intersection></hsegment></shape></wire>
<wire>
<ID>784 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-204,90.5,-204</points>
<connection>
<GID>545</GID>
<name>IN_0</name></connection>
<connection>
<GID>534</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>767 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-176.5,245.5,-176.5</points>
<connection>
<GID>513</GID>
<name>IN_0</name></connection>
<connection>
<GID>510</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>954 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-178.5,245.5,-178.5</points>
<connection>
<GID>513</GID>
<name>IN_1</name></connection>
<connection>
<GID>710</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>773 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,-177.5,270.5,-162.5</points>
<intersection>-177.5 2</intersection>
<intersection>-162.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>251.5,-177.5,270.5,-177.5</points>
<connection>
<GID>513</GID>
<name>OUT</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>270.5,-162.5,271,-162.5</points>
<connection>
<GID>529</GID>
<name>IN_5</name></connection>
<intersection>270.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>756 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-146.5,245.5,-146.5</points>
<connection>
<GID>517</GID>
<name>IN_0</name></connection>
<connection>
<GID>507</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>760 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-158.5,245.5,-158.5</points>
<connection>
<GID>521</GID>
<name>IN_0</name></connection>
<connection>
<GID>509</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>896 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-121.5,87,-121.5</points>
<connection>
<GID>344</GID>
<name>IN_0</name></connection>
<connection>
<GID>649</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>927 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-160.5,90.5,-160.5</points>
<connection>
<GID>680</GID>
<name>IN_0</name></connection>
<connection>
<GID>434</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>952 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>241.5,-166.5,241.5,-166.5</points>
<connection>
<GID>525</GID>
<name>IN_0</name></connection>
<connection>
<GID>708</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>630 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167,-126.5,167,-116.5</points>
<intersection>-126.5 2</intersection>
<intersection>-116.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>167,-116.5,168,-116.5</points>
<connection>
<GID>376</GID>
<name>IN_6</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148.5,-126.5,167,-126.5</points>
<connection>
<GID>359</GID>
<name>OUT</name></connection>
<intersection>167 0</intersection></hsegment></shape></wire>
<wire>
<ID>989 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123.5,-115,123.5,-115</points>
<connection>
<GID>349</GID>
<name>OUT</name></connection>
<connection>
<GID>745</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>745 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219.5,-156.5,219.5,-140.5</points>
<connection>
<GID>504</GID>
<name>IN_0</name></connection>
<intersection>-140.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>200,-140.5,219.5,-140.5</points>
<connection>
<GID>483</GID>
<name>OUT</name></connection>
<intersection>219.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>770 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,-157.5,270.5,-147.5</points>
<intersection>-157.5 1</intersection>
<intersection>-147.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>270.5,-157.5,271,-157.5</points>
<connection>
<GID>529</GID>
<name>IN_1</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>251.5,-147.5,270.5,-147.5</points>
<connection>
<GID>507</GID>
<name>OUT</name></connection>
<intersection>270.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>771 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270,-158.5,270,-153.5</points>
<intersection>-158.5 1</intersection>
<intersection>-153.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>270,-158.5,271,-158.5</points>
<connection>
<GID>529</GID>
<name>IN_2</name></connection>
<intersection>270 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>251.5,-153.5,270,-153.5</points>
<connection>
<GID>508</GID>
<name>OUT</name></connection>
<intersection>270 0</intersection></hsegment></shape></wire>
<wire>
<ID>649 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>220,-111.5,220,-95.5</points>
<connection>
<GID>399</GID>
<name>IN_0</name></connection>
<intersection>-95.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>200.5,-95.5,220,-95.5</points>
<connection>
<GID>378</GID>
<name>OUT</name></connection>
<intersection>220 0</intersection></hsegment></shape></wire>
<wire>
<ID>472 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271,-164,271,-163.5</points>
<connection>
<GID>529</GID>
<name>IN_4</name></connection>
<connection>
<GID>224</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>996 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278,-160,278,-160</points>
<connection>
<GID>529</GID>
<name>OUT</name></connection>
<connection>
<GID>752</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>609 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-93.5,142.5,-93.5</points>
<connection>
<GID>352</GID>
<name>IN_0</name></connection>
<connection>
<GID>361</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>899 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-95.5,142.5,-95.5</points>
<connection>
<GID>352</GID>
<name>IN_1</name></connection>
<connection>
<GID>652</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>900 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-97.5,142.5,-97.5</points>
<connection>
<GID>352</GID>
<name>IN_2</name></connection>
<connection>
<GID>653</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>625 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168,-111.5,168,-95.5</points>
<connection>
<GID>376</GID>
<name>IN_0</name></connection>
<intersection>-95.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>148.5,-95.5,168,-95.5</points>
<connection>
<GID>352</GID>
<name>OUT</name></connection>
<intersection>168 0</intersection></hsegment></shape></wire>
<wire>
<ID>933 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-148.5,142,-148.5</points>
<connection>
<GID>688</GID>
<name>IN_0</name></connection>
<connection>
<GID>458</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>985 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-224,245.5,-224</points>
<connection>
<GID>609</GID>
<name>IN_1</name></connection>
<connection>
<GID>741</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>626 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167.5,-112.5,167.5,-102.5</points>
<intersection>-112.5 1</intersection>
<intersection>-102.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>167.5,-112.5,168,-112.5</points>
<connection>
<GID>376</GID>
<name>IN_1</name></connection>
<intersection>167.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148.5,-102.5,167.5,-102.5</points>
<connection>
<GID>353</GID>
<name>OUT</name></connection>
<intersection>167.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>997 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,-205.5,123,-205.5</points>
<connection>
<GID>554</GID>
<name>OUT</name></connection>
<connection>
<GID>753</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>638 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-107.5,194.5,-107.5</points>
<connection>
<GID>354</GID>
<name>IN_0</name></connection>
<connection>
<GID>388</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>910 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-109.5,194.5,-109.5</points>
<connection>
<GID>354</GID>
<name>IN_1</name></connection>
<connection>
<GID>663</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>651 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219,-113.5,219,-108.5</points>
<intersection>-113.5 1</intersection>
<intersection>-108.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>219,-113.5,220,-113.5</points>
<connection>
<GID>399</GID>
<name>IN_2</name></connection>
<intersection>219 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200.5,-108.5,219,-108.5</points>
<connection>
<GID>354</GID>
<name>OUT</name></connection>
<intersection>219 0</intersection></hsegment></shape></wire>
<wire>
<ID>962 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-224,90.5,-224</points>
<connection>
<GID>718</GID>
<name>IN_0</name></connection>
<connection>
<GID>537</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>973 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-194,194,-194</points>
<connection>
<GID>583</GID>
<name>IN_1</name></connection>
<connection>
<GID>729</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>614 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-107.5,142.5,-107.5</points>
<connection>
<GID>355</GID>
<name>IN_0</name></connection>
<connection>
<GID>366</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>902 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-109.5,142.5,-109.5</points>
<connection>
<GID>355</GID>
<name>IN_1</name></connection>
<connection>
<GID>655</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>958 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-200,90.5,-200</points>
<connection>
<GID>533</GID>
<name>IN_1</name></connection>
<connection>
<GID>714</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>795 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-204,115,-199</points>
<intersection>-204 1</intersection>
<intersection>-199 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,-204,116,-204</points>
<connection>
<GID>554</GID>
<name>IN_2</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>96.5,-199,115,-199</points>
<connection>
<GID>533</GID>
<name>OUT</name></connection>
<intersection>115 0</intersection></hsegment></shape></wire>
<wire>
<ID>937 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-172.5,142,-172.5</points>
<connection>
<GID>692</GID>
<name>IN_0</name></connection>
<connection>
<GID>464</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>977 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-218,194,-218</points>
<connection>
<GID>585</GID>
<name>IN_1</name></connection>
<connection>
<GID>733</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>618 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-119.5,142.5,-119.5</points>
<connection>
<GID>358</GID>
<name>IN_0</name></connection>
<connection>
<GID>370</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>950 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-154.5,245.5,-154.5</points>
<connection>
<GID>706</GID>
<name>IN_0</name></connection>
<connection>
<GID>508</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>791 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-222,90.5,-222</points>
<connection>
<GID>537</GID>
<name>IN_0</name></connection>
<connection>
<GID>552</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>906 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-133.5,142.5,-133.5</points>
<connection>
<GID>360</GID>
<name>IN_1</name></connection>
<connection>
<GID>659</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>629 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167.5,-132.5,167.5,-117.5</points>
<intersection>-132.5 2</intersection>
<intersection>-117.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>148.5,-132.5,167.5,-132.5</points>
<connection>
<GID>360</GID>
<name>OUT</name></connection>
<intersection>167.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>167.5,-117.5,168,-117.5</points>
<connection>
<GID>376</GID>
<name>IN_5</name></connection>
<intersection>167.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>941 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-148.5,194,-148.5</points>
<connection>
<GID>696</GID>
<name>IN_0</name></connection>
<connection>
<GID>484</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>960 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,-212,86.5,-212</points>
<connection>
<GID>549</GID>
<name>IN_0</name></connection>
<connection>
<GID>716</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>787 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-212,90.5,-212</points>
<connection>
<GID>549</GID>
<name>OUT_0</name></connection>
<connection>
<GID>535</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>904 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,-121.5,138.5,-121.5</points>
<connection>
<GID>372</GID>
<name>IN_0</name></connection>
<connection>
<GID>657</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>819 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166.5,-204,166.5,-199</points>
<intersection>-204 1</intersection>
<intersection>-199 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166.5,-204,167.5,-204</points>
<connection>
<GID>580</GID>
<name>IN_2</name></connection>
<intersection>166.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148,-199,166.5,-199</points>
<connection>
<GID>560</GID>
<name>OUT</name></connection>
<intersection>166.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>322 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167.5,-209.5,167.5,-209</points>
<connection>
<GID>580</GID>
<name>IN_4</name></connection>
<connection>
<GID>152</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>823 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,-211,166,-206</points>
<intersection>-211 2</intersection>
<intersection>-206 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166,-206,167.5,-206</points>
<connection>
<GID>580</GID>
<name>IN_7</name></connection>
<intersection>166 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148,-211,166,-211</points>
<connection>
<GID>563</GID>
<name>OUT</name></connection>
<intersection>166 0</intersection></hsegment></shape></wire>
<wire>
<ID>681 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-138.5,90.5,-138.5</points>
<connection>
<GID>430</GID>
<name>IN_0</name></connection>
<connection>
<GID>438</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>504 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168,-119,168,-118.5</points>
<connection>
<GID>376</GID>
<name>IN_4</name></connection>
<connection>
<GID>229</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>834 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-210,194,-210</points>
<connection>
<GID>584</GID>
<name>IN_0</name></connection>
<connection>
<GID>593</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>835 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-212,194,-212</points>
<connection>
<GID>584</GID>
<name>IN_1</name></connection>
<connection>
<GID>595</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>486 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271.5,-119,271.5,-118.5</points>
<connection>
<GID>424</GID>
<name>IN_4</name></connection>
<connection>
<GID>225</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>328 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116,-164,116,-163.5</points>
<connection>
<GID>454</GID>
<name>IN_4</name></connection>
<connection>
<GID>164</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>633 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-93.5,194.5,-93.5</points>
<connection>
<GID>378</GID>
<name>IN_0</name></connection>
<connection>
<GID>384</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>908 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-97.5,194.5,-97.5</points>
<connection>
<GID>378</GID>
<name>IN_2</name></connection>
<connection>
<GID>661</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>650 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219.5,-112.5,219.5,-102.5</points>
<intersection>-112.5 1</intersection>
<intersection>-102.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>219.5,-112.5,220,-112.5</points>
<connection>
<GID>399</GID>
<name>IN_1</name></connection>
<intersection>219.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200.5,-102.5,219.5,-102.5</points>
<connection>
<GID>379</GID>
<name>OUT</name></connection>
<intersection>219.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>655 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218.5,-120.5,218.5,-115.5</points>
<intersection>-120.5 2</intersection>
<intersection>-115.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218.5,-115.5,220,-115.5</points>
<connection>
<GID>399</GID>
<name>IN_7</name></connection>
<intersection>218.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200.5,-120.5,218.5,-120.5</points>
<connection>
<GID>381</GID>
<name>OUT</name></connection>
<intersection>218.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>974 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-200,194,-200</points>
<connection>
<GID>730</GID>
<name>IN_0</name></connection>
<connection>
<GID>559</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>647 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-131.5,194.5,-131.5</points>
<connection>
<GID>383</GID>
<name>IN_0</name></connection>
<connection>
<GID>397</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>914 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-133.5,194.5,-133.5</points>
<connection>
<GID>383</GID>
<name>IN_1</name></connection>
<connection>
<GID>667</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>934 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-154.5,142,-154.5</points>
<connection>
<GID>689</GID>
<name>IN_0</name></connection>
<connection>
<GID>460</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>912 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190.5,-121.5,190.5,-121.5</points>
<connection>
<GID>394</GID>
<name>IN_0</name></connection>
<connection>
<GID>665</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>976 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190,-212,190,-212</points>
<connection>
<GID>732</GID>
<name>IN_0</name></connection>
<connection>
<GID>595</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>968 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-212,138,-212</points>
<connection>
<GID>577</GID>
<name>IN_0</name></connection>
<connection>
<GID>724</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>811 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-212,142,-212</points>
<connection>
<GID>577</GID>
<name>OUT_0</name></connection>
<connection>
<GID>563</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>660 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-101.5,246,-101.5</points>
<connection>
<GID>402</GID>
<name>IN_0</name></connection>
<connection>
<GID>412</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>674 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271,-112.5,271,-102.5</points>
<intersection>-112.5 1</intersection>
<intersection>-102.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>271,-112.5,271.5,-112.5</points>
<connection>
<GID>424</GID>
<name>IN_1</name></connection>
<intersection>271 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>252,-102.5,271,-102.5</points>
<connection>
<GID>402</GID>
<name>OUT</name></connection>
<intersection>271 0</intersection></hsegment></shape></wire>
<wire>
<ID>918 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-109.5,246,-109.5</points>
<connection>
<GID>403</GID>
<name>IN_1</name></connection>
<connection>
<GID>671</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>675 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,-113.5,270.5,-108.5</points>
<intersection>-113.5 1</intersection>
<intersection>-108.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>270.5,-113.5,271.5,-113.5</points>
<connection>
<GID>424</GID>
<name>IN_2</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>252,-108.5,270.5,-108.5</points>
<connection>
<GID>403</GID>
<name>OUT</name></connection>
<intersection>270.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>664 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-113.5,246,-113.5</points>
<connection>
<GID>404</GID>
<name>IN_0</name></connection>
<connection>
<GID>416</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>919 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-115.5,246,-115.5</points>
<connection>
<GID>404</GID>
<name>IN_1</name></connection>
<connection>
<GID>672</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>676 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>252,-114.5,271.5,-114.5</points>
<connection>
<GID>404</GID>
<name>OUT</name></connection>
<connection>
<GID>424</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>671 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-131.5,246,-131.5</points>
<connection>
<GID>405</GID>
<name>IN_0</name></connection>
<connection>
<GID>408</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>666 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-119.5,246,-119.5</points>
<connection>
<GID>406</GID>
<name>IN_0</name></connection>
<connection>
<GID>418</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>828 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-192,194,-192</points>
<connection>
<GID>589</GID>
<name>IN_0</name></connection>
<connection>
<GID>583</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>667 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-121.5,246,-121.5</points>
<connection>
<GID>406</GID>
<name>IN_1</name></connection>
<connection>
<GID>420</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>679 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270,-120.5,270,-115.5</points>
<intersection>-120.5 2</intersection>
<intersection>-115.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>270,-115.5,271.5,-115.5</points>
<connection>
<GID>424</GID>
<name>IN_7</name></connection>
<intersection>270 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>252,-120.5,270,-120.5</points>
<connection>
<GID>406</GID>
<name>OUT</name></connection>
<intersection>270 0</intersection></hsegment></shape></wire>
<wire>
<ID>921 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-127.5,246,-127.5</points>
<connection>
<GID>407</GID>
<name>IN_1</name></connection>
<connection>
<GID>674</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>678 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,-126.5,270.5,-116.5</points>
<intersection>-126.5 2</intersection>
<intersection>-116.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>270.5,-116.5,271.5,-116.5</points>
<connection>
<GID>424</GID>
<name>IN_6</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>252,-126.5,270.5,-126.5</points>
<connection>
<GID>407</GID>
<name>OUT</name></connection>
<intersection>270.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>922 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,-133.5,246,-133.5</points>
<connection>
<GID>408</GID>
<name>IN_1</name></connection>
<connection>
<GID>675</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>923 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-140.5,90.5,-140.5</points>
<connection>
<GID>430</GID>
<name>IN_1</name></connection>
<connection>
<GID>676</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>697 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116,-156.5,116,-140.5</points>
<connection>
<GID>454</GID>
<name>IN_0</name></connection>
<intersection>-140.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>96.5,-140.5,116,-140.5</points>
<connection>
<GID>430</GID>
<name>OUT</name></connection>
<intersection>116 0</intersection></hsegment></shape></wire>
<wire>
<ID>863 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-222,245.5,-222</points>
<connection>
<GID>609</GID>
<name>IN_0</name></connection>
<connection>
<GID>606</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>684 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-146.5,90.5,-146.5</points>
<connection>
<GID>432</GID>
<name>IN_0</name></connection>
<connection>
<GID>441</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>698 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-157.5,115.5,-147.5</points>
<intersection>-157.5 1</intersection>
<intersection>-147.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115.5,-157.5,116,-157.5</points>
<connection>
<GID>454</GID>
<name>IN_1</name></connection>
<intersection>115.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>96.5,-147.5,115.5,-147.5</points>
<connection>
<GID>432</GID>
<name>OUT</name></connection>
<intersection>115.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>686 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-152.5,90.5,-152.5</points>
<connection>
<GID>433</GID>
<name>IN_0</name></connection>
<connection>
<GID>443</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>926 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-154.5,90.5,-154.5</points>
<connection>
<GID>433</GID>
<name>IN_1</name></connection>
<connection>
<GID>679</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>699 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-158.5,115,-153.5</points>
<intersection>-158.5 1</intersection>
<intersection>-153.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,-158.5,116,-158.5</points>
<connection>
<GID>454</GID>
<name>IN_2</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>96.5,-153.5,115,-153.5</points>
<connection>
<GID>433</GID>
<name>OUT</name></connection>
<intersection>115 0</intersection></hsegment></shape></wire>
<wire>
<ID>688 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-158.5,90.5,-158.5</points>
<connection>
<GID>434</GID>
<name>IN_0</name></connection>
<connection>
<GID>445</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>700 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96.5,-159.5,116,-159.5</points>
<connection>
<GID>434</GID>
<name>OUT</name></connection>
<connection>
<GID>454</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>690 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-164.5,90.5,-164.5</points>
<connection>
<GID>435</GID>
<name>IN_0</name></connection>
<connection>
<GID>447</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>691 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-166.5,90.5,-166.5</points>
<connection>
<GID>435</GID>
<name>IN_1</name></connection>
<connection>
<GID>449</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>703 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-165.5,114.5,-160.5</points>
<intersection>-165.5 2</intersection>
<intersection>-160.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,-160.5,116,-160.5</points>
<connection>
<GID>454</GID>
<name>IN_7</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>96.5,-165.5,114.5,-165.5</points>
<connection>
<GID>435</GID>
<name>OUT</name></connection>
<intersection>114.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>852 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-192,245.5,-192</points>
<connection>
<GID>613</GID>
<name>IN_0</name></connection>
<connection>
<GID>603</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>693 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-170.5,90.5,-170.5</points>
<connection>
<GID>436</GID>
<name>IN_0</name></connection>
<connection>
<GID>450</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>702 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-171.5,115,-161.5</points>
<intersection>-171.5 2</intersection>
<intersection>-161.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,-161.5,116,-161.5</points>
<connection>
<GID>454</GID>
<name>IN_6</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>96.5,-171.5,115,-171.5</points>
<connection>
<GID>436</GID>
<name>OUT</name></connection>
<intersection>115 0</intersection></hsegment></shape></wire>
<wire>
<ID>695 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-176.5,90.5,-176.5</points>
<connection>
<GID>437</GID>
<name>IN_0</name></connection>
<connection>
<GID>452</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>930 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-178.5,90.5,-178.5</points>
<connection>
<GID>437</GID>
<name>IN_1</name></connection>
<connection>
<GID>683</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>701 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-177.5,115.5,-162.5</points>
<intersection>-177.5 2</intersection>
<intersection>-162.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>96.5,-177.5,115.5,-177.5</points>
<connection>
<GID>437</GID>
<name>OUT</name></connection>
<intersection>115.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>115.5,-162.5,116,-162.5</points>
<connection>
<GID>454</GID>
<name>IN_5</name></connection>
<intersection>115.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>928 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,-166.5,86.5,-166.5</points>
<connection>
<GID>449</GID>
<name>IN_0</name></connection>
<connection>
<GID>681</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>981 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-194,245.5,-194</points>
<connection>
<GID>603</GID>
<name>IN_1</name></connection>
<connection>
<GID>737</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>993 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,-160,123,-160</points>
<connection>
<GID>454</GID>
<name>OUT</name></connection>
<connection>
<GID>749</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>858 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-210,245.5,-210</points>
<connection>
<GID>607</GID>
<name>IN_0</name></connection>
<connection>
<GID>618</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>705 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-138.5,142,-138.5</points>
<connection>
<GID>457</GID>
<name>IN_0</name></connection>
<connection>
<GID>466</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>931 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-140.5,142,-140.5</points>
<connection>
<GID>457</GID>
<name>IN_1</name></connection>
<connection>
<GID>686</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>932 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-142.5,142,-142.5</points>
<connection>
<GID>457</GID>
<name>IN_2</name></connection>
<connection>
<GID>687</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>758 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-152.5,245.5,-152.5</points>
<connection>
<GID>519</GID>
<name>IN_0</name></connection>
<connection>
<GID>508</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>939 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-140.5,194,-140.5</points>
<connection>
<GID>483</GID>
<name>IN_1</name></connection>
<connection>
<GID>694</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>940 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-142.5,194,-142.5</points>
<connection>
<GID>483</GID>
<name>IN_2</name></connection>
<connection>
<GID>695</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>732 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-146.5,194,-146.5</points>
<connection>
<GID>484</GID>
<name>IN_0</name></connection>
<connection>
<GID>491</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>746 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219,-157.5,219,-147.5</points>
<intersection>-157.5 1</intersection>
<intersection>-147.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>219,-157.5,219.5,-157.5</points>
<connection>
<GID>504</GID>
<name>IN_1</name></connection>
<intersection>219 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200,-147.5,219,-147.5</points>
<connection>
<GID>484</GID>
<name>OUT</name></connection>
<intersection>219 0</intersection></hsegment></shape></wire>
<wire>
<ID>738 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-164.5,194,-164.5</points>
<connection>
<GID>486</GID>
<name>IN_0</name></connection>
<connection>
<GID>497</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>751 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>218,-165.5,218,-160.5</points>
<intersection>-165.5 2</intersection>
<intersection>-160.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>218,-160.5,219.5,-160.5</points>
<connection>
<GID>504</GID>
<name>IN_7</name></connection>
<intersection>218 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>200,-165.5,218,-165.5</points>
<connection>
<GID>486</GID>
<name>OUT</name></connection>
<intersection>218 0</intersection></hsegment></shape></wire>
<wire>
<ID>946 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-178.5,194,-178.5</points>
<connection>
<GID>488</GID>
<name>IN_1</name></connection>
<connection>
<GID>702</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>948 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-142.5,245.5,-142.5</points>
<connection>
<GID>704</GID>
<name>IN_0</name></connection>
<connection>
<GID>506</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>799 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-211,114.5,-206</points>
<intersection>-211 2</intersection>
<intersection>-206 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,-206,116,-206</points>
<connection>
<GID>554</GID>
<name>IN_7</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>96.5,-211,114.5,-211</points>
<connection>
<GID>535</GID>
<name>OUT</name></connection>
<intersection>114.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>956 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-188,90.5,-188</points>
<connection>
<GID>712</GID>
<name>IN_0</name></connection>
<connection>
<GID>531</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>947 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-140.5,245.5,-140.5</points>
<connection>
<GID>506</GID>
<name>IN_1</name></connection>
<connection>
<GID>703</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>949 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-148.5,245.5,-148.5</points>
<connection>
<GID>507</GID>
<name>IN_1</name></connection>
<connection>
<GID>705</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>951 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-160.5,245.5,-160.5</points>
<connection>
<GID>509</GID>
<name>IN_1</name></connection>
<connection>
<GID>707</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>957 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-194,90.5,-194</points>
<connection>
<GID>532</GID>
<name>IN_1</name></connection>
<connection>
<GID>713</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>959 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-206,90.5,-206</points>
<connection>
<GID>534</GID>
<name>IN_1</name></connection>
<connection>
<GID>715</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>323 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116,-209.5,116,-209</points>
<connection>
<GID>554</GID>
<name>IN_4</name></connection>
<connection>
<GID>156</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>966 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-200,142,-200</points>
<connection>
<GID>560</GID>
<name>IN_1</name></connection>
<connection>
<GID>722</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>969 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-218,142,-218</points>
<connection>
<GID>564</GID>
<name>IN_1</name></connection>
<connection>
<GID>725</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>972 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-188,194,-188</points>
<connection>
<GID>582</GID>
<name>IN_2</name></connection>
<connection>
<GID>728</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>839 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-222,194,-222</points>
<connection>
<GID>586</GID>
<name>IN_0</name></connection>
<connection>
<GID>598</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>978 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-224,194,-224</points>
<connection>
<GID>586</GID>
<name>IN_1</name></connection>
<connection>
<GID>734</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>849 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-184,245.5,-184</points>
<connection>
<GID>602</GID>
<name>IN_0</name></connection>
<connection>
<GID>610</GID>
<name>IN_0</name></connection></vsegment></shape></wire></page 1>
<page 2>
<PageViewport>-199.633,28.894,389.305,-263.465</PageViewport>
<gate>
<ID>315</ID>
<type>DA_FROM</type>
<position>96.5,-19</position>
<input>
<ID>IN_0</ID>615 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>1024</ID>
<type>AA_LABEL</type>
<position>37.5,-32.5</position>
<gparam>LABEL_TEXT E Set/Reset</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>845</ID>
<type>AE_OR2</type>
<position>189,-85</position>
<input>
<ID>IN_0</ID>345 </input>
<input>
<ID>IN_1</ID>1045 </input>
<output>
<ID>OUT</ID>1043 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>140</ID>
<type>AA_AND2</type>
<position>249.5,-24.5</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>150 </input>
<output>
<ID>OUT</ID>584 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>957</ID>
<type>DA_FROM</type>
<position>217.5,-31.5</position>
<input>
<ID>IN_0</ID>1122 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>389</ID>
<type>BE_DECODER_3x8</type>
<position>-109,-24</position>
<input>
<ID>ENABLE</ID>692 </input>
<input>
<ID>IN_0</ID>661 </input>
<input>
<ID>IN_1</ID>663 </input>
<input>
<ID>IN_2</ID>665 </input>
<output>
<ID>OUT_0</ID>680 </output>
<output>
<ID>OUT_1</ID>687 </output>
<output>
<ID>OUT_2</ID>670 </output>
<output>
<ID>OUT_3</ID>685 </output>
<output>
<ID>OUT_4</ID>668 </output>
<output>
<ID>OUT_5</ID>683 </output>
<output>
<ID>OUT_6</ID>672 </output>
<output>
<ID>OUT_7</ID>682 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>883</ID>
<type>AE_SMALL_INVERTER</type>
<position>143.5,-172</position>
<input>
<ID>IN_0</ID>1074 </input>
<output>
<ID>OUT_0</ID>1076 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1247</ID>
<type>DE_TO</type>
<position>-38,-114</position>
<input>
<ID>IN_0</ID>1360 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHL</lparam></gate>
<gate>
<ID>396</ID>
<type>DA_FROM</type>
<position>-114,-25.5</position>
<input>
<ID>IN_0</ID>665 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir14</lparam></gate>
<gate>
<ID>617</ID>
<type>AA_LABEL</type>
<position>131.5,-71.5</position>
<gparam>LABEL_TEXT PC Commands</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>440</ID>
<type>AA_LABEL</type>
<position>-107.5,-15</position>
<gparam>LABEL_TEXT Instruction Decoder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>553</ID>
<type>AE_OR2</type>
<position>100,-56</position>
<input>
<ID>IN_0</ID>759 </input>
<input>
<ID>IN_1</ID>761 </input>
<output>
<ID>OUT</ID>757 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>448</ID>
<type>DA_FROM</type>
<position>148.5,-16</position>
<input>
<ID>IN_0</ID>711 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>468</ID>
<type>DA_FROM</type>
<position>142.5,-25</position>
<input>
<ID>IN_0</ID>709 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>1241</ID>
<type>DE_TO</type>
<position>-38,-80.5</position>
<input>
<ID>IN_0</ID>1340 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>398</ID>
<type>DE_TO</type>
<position>-104,-25.5</position>
<input>
<ID>IN_0</ID>670 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>334</ID>
<type>DA_FROM</type>
<position>100.5,-23</position>
<input>
<ID>IN_0</ID>641 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T3</lparam></gate>
<gate>
<ID>245</ID>
<type>DA_FROM</type>
<position>16,-69</position>
<input>
<ID>IN_0</ID>350 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B10</lparam></gate>
<gate>
<ID>1113</ID>
<type>DA_FROM</type>
<position>27.5,-114.5</position>
<input>
<ID>IN_0</ID>1237 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>964</ID>
<type>DE_TO</type>
<position>230.5,-22.5</position>
<input>
<ID>IN_0</ID>1131 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>249</ID>
<type>AE_OR4</type>
<position>34.5,-62</position>
<input>
<ID>IN_0</ID>352 </input>
<input>
<ID>IN_1</ID>353 </input>
<input>
<ID>IN_2</ID>354 </input>
<input>
<ID>IN_3</ID>355 </input>
<output>
<ID>OUT</ID>351 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>968</ID>
<type>AA_REGISTER4</type>
<position>218.5,-25.5</position>
<output>
<ID>OUT_0</ID>1125 </output>
<output>
<ID>OUT_1</ID>1126 </output>
<output>
<ID>OUT_2</ID>1124 </output>
<input>
<ID>clear</ID>1136 </input>
<input>
<ID>clock</ID>1122 </input>
<input>
<ID>count_enable</ID>600 </input>
<input>
<ID>count_up</ID>600 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>805</ID>
<type>AA_AND2</type>
<position>142.5,-106</position>
<input>
<ID>IN_0</ID>1005 </input>
<input>
<ID>IN_1</ID>1004 </input>
<output>
<ID>OUT</ID>1034 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>467</ID>
<type>DA_FROM</type>
<position>142.5,-23</position>
<input>
<ID>IN_0</ID>706 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>275</ID>
<type>DM_NOR8</type>
<position>-43.5,-37.5</position>
<input>
<ID>IN_0</ID>357 </input>
<input>
<ID>IN_1</ID>360 </input>
<input>
<ID>IN_2</ID>358 </input>
<input>
<ID>IN_3</ID>361 </input>
<input>
<ID>IN_4</ID>363 </input>
<input>
<ID>IN_5</ID>359 </input>
<input>
<ID>IN_6</ID>362 </input>
<input>
<ID>IN_7</ID>356 </input>
<output>
<ID>OUT</ID>380 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>766</ID>
<type>AE_SMALL_INVERTER</type>
<position>137.5,-81.5</position>
<input>
<ID>IN_0</ID>831 </input>
<output>
<ID>OUT_0</ID>1022 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1281</ID>
<type>DA_FROM</type>
<position>-44.5,-138</position>
<input>
<ID>IN_0</ID>1366 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir5</lparam></gate>
<gate>
<ID>413</ID>
<type>DE_TO</type>
<position>-104,-23.5</position>
<input>
<ID>IN_0</ID>668 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>285</ID>
<type>CC_PULSE</type>
<position>255,-21.5</position>
<output>
<ID>OUT_0</ID>560 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 40</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>971</ID>
<type>EE_VDD</type>
<position>222.5,-17.5</position>
<output>
<ID>OUT_0</ID>1135 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1110</ID>
<type>DA_FROM</type>
<position>27.5,-112.5</position>
<input>
<ID>IN_0</ID>1234 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B6</lparam></gate>
<gate>
<ID>417</ID>
<type>DE_TO</type>
<position>-104,-21.5</position>
<input>
<ID>IN_0</ID>672 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>991</ID>
<type>DA_FROM</type>
<position>228.5,-51.5</position>
<input>
<ID>IN_0</ID>1140 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>289</ID>
<type>DE_TO</type>
<position>116.5,-21</position>
<input>
<ID>IN_0</ID>646 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mem_read</lparam></gate>
<gate>
<ID>296</ID>
<type>DA_FROM</type>
<position>96.5,-13</position>
<input>
<ID>IN_0</ID>613 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>1151</ID>
<type>DA_FROM</type>
<position>49,-130</position>
<input>
<ID>IN_0</ID>1266 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>300</ID>
<type>AE_SMALL_INVERTER</type>
<position>100.5,-13</position>
<input>
<ID>IN_0</ID>613 </input>
<output>
<ID>OUT_0</ID>637 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1188</ID>
<type>AA_AND2</type>
<position>-36.5,-41.5</position>
<input>
<ID>IN_0</ID>380 </input>
<input>
<ID>IN_1</ID>389 </input>
<output>
<ID>OUT</ID>1296 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>503</ID>
<type>AA_LABEL</type>
<position>132,-40.5</position>
<gparam>LABEL_TEXT AR Commands</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>311</ID>
<type>DA_FROM</type>
<position>100.5,-15</position>
<input>
<ID>IN_0</ID>635 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T1</lparam></gate>
<gate>
<ID>319</ID>
<type>AE_SMALL_INVERTER</type>
<position>100.5,-19</position>
<input>
<ID>IN_0</ID>615 </input>
<output>
<ID>OUT_0</ID>644 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>789</ID>
<type>DA_FROM</type>
<position>125.5,-123.5</position>
<input>
<ID>IN_0</ID>1012 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B9</lparam></gate>
<gate>
<ID>451</ID>
<type>DA_FROM</type>
<position>148.5,-18</position>
<input>
<ID>IN_0</ID>713 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T1</lparam></gate>
<gate>
<ID>387</ID>
<type>AE_OR3</type>
<position>111.5,-21</position>
<input>
<ID>IN_0</ID>648 </input>
<input>
<ID>IN_1</ID>658 </input>
<input>
<ID>IN_2</ID>659 </input>
<output>
<ID>OUT</ID>646 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>323</ID>
<type>DA_FROM</type>
<position>100.5,-21</position>
<input>
<ID>IN_0</ID>639 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID I</lparam></gate>
<gate>
<ID>1030</ID>
<type>DA_FROM</type>
<position>16,-44</position>
<input>
<ID>IN_0</ID>1169 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B6</lparam></gate>
<gate>
<ID>337</ID>
<type>DA_FROM</type>
<position>87.5,-25.5</position>
<input>
<ID>IN_0</ID>617 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>1028</ID>
<type>DA_FROM</type>
<position>16,-38</position>
<input>
<ID>IN_0</ID>1166 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>343</ID>
<type>DA_FROM</type>
<position>87.5,-27.5</position>
<input>
<ID>IN_0</ID>620 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>806</ID>
<type>AA_AND2</type>
<position>128.5,-114</position>
<input>
<ID>IN_0</ID>1010 </input>
<input>
<ID>IN_1</ID>1011 </input>
<output>
<ID>OUT</ID>1009 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>476</ID>
<type>AE_OR2</type>
<position>147.5,-22</position>
<input>
<ID>IN_0</ID>704 </input>
<input>
<ID>IN_1</ID>706 </input>
<output>
<ID>OUT</ID>707 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1199</ID>
<type>DA_FROM</type>
<position>-56,-39</position>
<input>
<ID>IN_0</ID>362 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr5</lparam></gate>
<gate>
<ID>348</ID>
<type>DA_FROM</type>
<position>87.5,-29.5</position>
<input>
<ID>IN_0</ID>622 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>1100</ID>
<type>AA_AND2</type>
<position>43.5,-92</position>
<input>
<ID>IN_0</ID>1225 </input>
<input>
<ID>IN_1</ID>1224 </input>
<output>
<ID>OUT</ID>1227 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>415</ID>
<type>DE_TO</type>
<position>-99,-22.5</position>
<input>
<ID>IN_0</ID>683 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>351</ID>
<type>DA_FROM</type>
<position>87.5,-31.5</position>
<input>
<ID>IN_0</ID>624 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>527</ID>
<type>DA_FROM</type>
<position>84.5,-59</position>
<input>
<ID>IN_0</ID>148 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>490</ID>
<type>AA_AND2</type>
<position>153.5,-17</position>
<input>
<ID>IN_0</ID>711 </input>
<input>
<ID>IN_1</ID>713 </input>
<output>
<ID>OUT</ID>730 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>426</ID>
<type>EE_VDD</type>
<position>-112,-18.5</position>
<output>
<ID>OUT_0</ID>692 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>362</ID>
<type>DA_FROM</type>
<position>87.5,-33.5</position>
<input>
<ID>IN_0</ID>634 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>365</ID>
<type>AE_OR4</type>
<position>98.5,-28.5</position>
<input>
<ID>IN_0</ID>617 </input>
<input>
<ID>IN_1</ID>620 </input>
<input>
<ID>IN_2</ID>622 </input>
<input>
<ID>IN_3</ID>624 </input>
<output>
<ID>OUT</ID>632 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1062</ID>
<type>DA_FROM</type>
<position>44.5,-87</position>
<input>
<ID>IN_0</ID>1197 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>576</ID>
<type>DA_FROM</type>
<position>141,-55</position>
<input>
<ID>IN_0</ID>778 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>369</ID>
<type>AA_AND2</type>
<position>105.5,-29.5</position>
<input>
<ID>IN_0</ID>632 </input>
<input>
<ID>IN_1</ID>634 </input>
<output>
<ID>OUT</ID>659 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>374</ID>
<type>AA_AND2</type>
<position>105.5,-14</position>
<input>
<ID>IN_0</ID>637 </input>
<input>
<ID>IN_1</ID>635 </input>
<output>
<ID>OUT</ID>648 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>BE_JKFF_LOW</type>
<position>267.5,-23.5</position>
<input>
<ID>J</ID>560 </input>
<input>
<ID>K</ID>586 </input>
<output>
<ID>Q</ID>96 </output>
<input>
<ID>clock</ID>343 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1198</ID>
<type>DA_FROM</type>
<position>-48.5,-38</position>
<input>
<ID>IN_0</ID>356 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr4</lparam></gate>
<gate>
<ID>505</ID>
<type>DE_TO</type>
<position>105,-56</position>
<input>
<ID>IN_0</ID>757 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ldAR</lparam></gate>
<gate>
<ID>1070</ID>
<type>AE_SMALL_INVERTER</type>
<position>24.5,-85.5</position>
<input>
<ID>IN_0</ID>1200 </input>
<output>
<ID>OUT_0</ID>1221 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>377</ID>
<type>AA_AND3</type>
<position>105.5,-21</position>
<input>
<ID>IN_0</ID>644 </input>
<input>
<ID>IN_1</ID>639 </input>
<input>
<ID>IN_2</ID>641 </input>
<output>
<ID>OUT</ID>658 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>455</ID>
<type>DA_FROM</type>
<position>142.5,-21</position>
<input>
<ID>IN_0</ID>704 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>1204</ID>
<type>DA_FROM</type>
<position>-48.5,-44</position>
<input>
<ID>IN_0</ID>381 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr10</lparam></gate>
<gate>
<ID>391</ID>
<type>DA_FROM</type>
<position>-114,-27.5</position>
<input>
<ID>IN_0</ID>661 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir12</lparam></gate>
<gate>
<ID>393</ID>
<type>DA_FROM</type>
<position>-120.5,-26.5</position>
<input>
<ID>IN_0</ID>663 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir13</lparam></gate>
<gate>
<ID>400</ID>
<type>DE_TO</type>
<position>-104,-27.5</position>
<input>
<ID>IN_0</ID>680 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>410</ID>
<type>DE_TO</type>
<position>-99,-26.5</position>
<input>
<ID>IN_0</ID>687 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>1295</ID>
<type>DE_TO</type>
<position>-40.5,-140</position>
<input>
<ID>IN_0</ID>1367 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B6</lparam></gate>
<gate>
<ID>411</ID>
<type>DE_TO</type>
<position>-99,-24.5</position>
<input>
<ID>IN_0</ID>685 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>419</ID>
<type>DE_TO</type>
<position>-99,-20.5</position>
<input>
<ID>IN_0</ID>682 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>444</ID>
<type>DE_TO</type>
<position>164.5,-23</position>
<input>
<ID>IN_0</ID>720 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID mem_write</lparam></gate>
<gate>
<ID>619</ID>
<type>DE_TO</type>
<position>90,-84.5</position>
<input>
<ID>IN_0</ID>816 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ldPC</lparam></gate>
<gate>
<ID>470</ID>
<type>DA_FROM</type>
<position>148.5,-29</position>
<input>
<ID>IN_0</ID>716 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T6</lparam></gate>
<gate>
<ID>472</ID>
<type>DA_FROM</type>
<position>148.5,-27</position>
<input>
<ID>IN_0</ID>718 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>810</ID>
<type>AA_AND2</type>
<position>130.5,-122.5</position>
<input>
<ID>IN_0</ID>1013 </input>
<input>
<ID>IN_1</ID>1012 </input>
<output>
<ID>OUT</ID>1028 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>480</ID>
<type>AA_AND2</type>
<position>153.5,-23</position>
<input>
<ID>IN_0</ID>707 </input>
<input>
<ID>IN_1</ID>709 </input>
<output>
<ID>OUT</ID>728 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>515</ID>
<type>DA_FROM</type>
<position>79,-49.5</position>
<input>
<ID>IN_0</ID>733 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>494</ID>
<type>AA_AND2</type>
<position>153.5,-28</position>
<input>
<ID>IN_0</ID>718 </input>
<input>
<ID>IN_1</ID>716 </input>
<output>
<ID>OUT</ID>731 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>498</ID>
<type>AE_OR3</type>
<position>159.5,-23</position>
<input>
<ID>IN_0</ID>730 </input>
<input>
<ID>IN_1</ID>728 </input>
<input>
<ID>IN_2</ID>731 </input>
<output>
<ID>OUT</ID>720 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>501</ID>
<type>AA_LABEL</type>
<position>128.5,-3</position>
<gparam>LABEL_TEXT Memory Commands</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>995</ID>
<type>DA_FROM</type>
<position>241.5,-69</position>
<input>
<ID>IN_0</ID>1158 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>516</ID>
<type>AE_SMALL_INVERTER</type>
<position>83,-49.5</position>
<input>
<ID>IN_0</ID>733 </input>
<output>
<ID>OUT_0</ID>744 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1005</ID>
<type>AA_AND2</type>
<position>240.5,-58</position>
<input>
<ID>IN_0</ID>1146 </input>
<input>
<ID>IN_1</ID>1147 </input>
<output>
<ID>OUT</ID>1155 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>518</ID>
<type>DA_FROM</type>
<position>83,-51.5</position>
<input>
<ID>IN_0</ID>740 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T0</lparam></gate>
<gate>
<ID>317</ID>
<type>AA_AND2</type>
<position>272,-36.5</position>
<input>
<ID>IN_0</ID>565 </input>
<input>
<ID>IN_1</ID>574 </input>
<output>
<ID>OUT</ID>563 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1003</ID>
<type>AE_OR2</type>
<position>234.5,-57</position>
<input>
<ID>IN_0</ID>1144 </input>
<input>
<ID>IN_1</ID>1145 </input>
<output>
<ID>OUT</ID>1146 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>524</ID>
<type>DA_FROM</type>
<position>83,-53.5</position>
<input>
<ID>IN_0</ID>737 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T2</lparam></gate>
<gate>
<ID>528</ID>
<type>DA_FROM</type>
<position>88.5,-63</position>
<input>
<ID>IN_0</ID>755 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T3</lparam></gate>
<gate>
<ID>1017</ID>
<type>DA_FROM</type>
<position>244.5,-25.5</position>
<input>
<ID>IN_0</ID>150 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B0</lparam></gate>
<gate>
<ID>530</ID>
<type>DA_FROM</type>
<position>88.5,-61</position>
<input>
<ID>IN_0</ID>754 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID I</lparam></gate>
<gate>
<ID>1226</ID>
<type>DA_FROM</type>
<position>-56,-54.5</position>
<input>
<ID>IN_0</ID>395 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac3</lparam></gate>
<gate>
<ID>1019</ID>
<type>DE_TO</type>
<position>61,-18.5</position>
<input>
<ID>IN_0</ID>1243 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID I</lparam></gate>
<gate>
<ID>540</ID>
<type>AE_OR2</type>
<position>88,-52.5</position>
<input>
<ID>IN_0</ID>740 </input>
<input>
<ID>IN_1</ID>737 </input>
<output>
<ID>OUT</ID>742 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>544</ID>
<type>AA_AND2</type>
<position>94,-51.5</position>
<input>
<ID>IN_0</ID>744 </input>
<input>
<ID>IN_1</ID>742 </input>
<output>
<ID>OUT</ID>759 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1234</ID>
<type>DA_FROM</type>
<position>-56,-62.5</position>
<input>
<ID>IN_0</ID>589 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac11</lparam></gate>
<gate>
<ID>899</ID>
<type>DE_TO</type>
<position>104,-214.5</position>
<input>
<ID>IN_0</ID>1103 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ldAC</lparam></gate>
<gate>
<ID>548</ID>
<type>AA_AND3</type>
<position>93.5,-61</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>754 </input>
<input>
<ID>IN_2</ID>755 </input>
<output>
<ID>OUT</ID>761 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>1249</ID>
<type>AA_AND2</type>
<position>-43,-80.5</position>
<input>
<ID>IN_0</ID>1341 </input>
<input>
<ID>IN_1</ID>1342 </input>
<output>
<ID>OUT</ID>1340 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>555</ID>
<type>DE_TO</type>
<position>127.5,-56</position>
<input>
<ID>IN_0</ID>776 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clrAR</lparam></gate>
<gate>
<ID>567</ID>
<type>DA_FROM</type>
<position>117.5,-55</position>
<input>
<ID>IN_0</ID>766 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>1285</ID>
<type>DA_FROM</type>
<position>-44.5,-146</position>
<input>
<ID>IN_0</ID>1370 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir9</lparam></gate>
<gate>
<ID>935</ID>
<type>AA_AND2</type>
<position>152.5,-215</position>
<input>
<ID>IN_0</ID>1107 </input>
<input>
<ID>IN_1</ID>1108 </input>
<output>
<ID>OUT</ID>1109 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>568</ID>
<type>DA_FROM</type>
<position>117.5,-57</position>
<input>
<ID>IN_0</ID>768 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T0</lparam></gate>
<gate>
<ID>1258</ID>
<type>AA_AND2</type>
<position>-43,-95</position>
<input>
<ID>IN_0</ID>1347 </input>
<input>
<ID>IN_1</ID>1348 </input>
<output>
<ID>OUT</ID>1349 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>572</ID>
<type>AA_AND2</type>
<position>122.5,-56</position>
<input>
<ID>IN_0</ID>766 </input>
<input>
<ID>IN_1</ID>768 </input>
<output>
<ID>OUT</ID>776 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1112</ID>
<type>AA_AND2</type>
<position>32.5,-111.5</position>
<input>
<ID>IN_0</ID>1233 </input>
<input>
<ID>IN_1</ID>1234 </input>
<output>
<ID>OUT</ID>1239 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>574</ID>
<type>DE_TO</type>
<position>151,-56</position>
<input>
<ID>IN_0</ID>781 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incAR</lparam></gate>
<gate>
<ID>579</ID>
<type>DA_FROM</type>
<position>141,-57</position>
<input>
<ID>IN_0</ID>779 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>1255</ID>
<type>DA_FROM</type>
<position>-48,-87</position>
<input>
<ID>IN_0</ID>1344 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>581</ID>
<type>AA_AND2</type>
<position>146,-56</position>
<input>
<ID>IN_0</ID>778 </input>
<input>
<ID>IN_1</ID>779 </input>
<output>
<ID>OUT</ID>781 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>588</ID>
<type>DE_TO</type>
<position>180.5,-56</position>
<input>
<ID>IN_0</ID>802 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID busAR</lparam></gate>
<gate>
<ID>1069</ID>
<type>AE_SMALL_INVERTER</type>
<position>24.5,-83.5</position>
<input>
<ID>IN_0</ID>1199 </input>
<output>
<ID>OUT_0</ID>1220 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>591</ID>
<type>DA_FROM</type>
<position>164,-53</position>
<input>
<ID>IN_0</ID>783 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>1283</ID>
<type>DA_FROM</type>
<position>-44.5,-142</position>
<input>
<ID>IN_0</ID>1368 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir7</lparam></gate>
<gate>
<ID>594</ID>
<type>DA_FROM</type>
<position>164,-55</position>
<input>
<ID>IN_0</ID>785 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>1271</ID>
<type>AA_AND2</type>
<position>-43,-114</position>
<input>
<ID>IN_0</ID>1358 </input>
<input>
<ID>IN_1</ID>1359 </input>
<output>
<ID>OUT</ID>1360 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>597</ID>
<type>AA_AND2</type>
<position>169,-54</position>
<input>
<ID>IN_0</ID>783 </input>
<input>
<ID>IN_1</ID>785 </input>
<output>
<ID>OUT</ID>792 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>599</ID>
<type>DA_FROM</type>
<position>164,-57</position>
<input>
<ID>IN_0</ID>788 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>601</ID>
<type>DA_FROM</type>
<position>164,-59</position>
<input>
<ID>IN_0</ID>790 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>611</ID>
<type>AA_AND2</type>
<position>169,-58</position>
<input>
<ID>IN_0</ID>788 </input>
<input>
<ID>IN_1</ID>790 </input>
<output>
<ID>OUT</ID>800 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>615</ID>
<type>AE_OR2</type>
<position>175.5,-56</position>
<input>
<ID>IN_0</ID>792 </input>
<input>
<ID>IN_1</ID>800 </input>
<output>
<ID>OUT</ID>802 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>623</ID>
<type>DA_FROM</type>
<position>73.5,-81.5</position>
<input>
<ID>IN_0</ID>803 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>625</ID>
<type>DA_FROM</type>
<position>73.5,-83.5</position>
<input>
<ID>IN_0</ID>805 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>626</ID>
<type>AA_AND2</type>
<position>78.5,-82.5</position>
<input>
<ID>IN_0</ID>803 </input>
<input>
<ID>IN_1</ID>805 </input>
<output>
<ID>OUT</ID>812 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>684</ID>
<type>DA_FROM</type>
<position>73.5,-85.5</position>
<input>
<ID>IN_0</ID>807 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>1231</ID>
<type>DA_FROM</type>
<position>-48.5,-59.5</position>
<input>
<ID>IN_0</ID>538 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac8</lparam></gate>
<gate>
<ID>685</ID>
<type>DA_FROM</type>
<position>73.5,-87.5</position>
<input>
<ID>IN_0</ID>809 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>697</ID>
<type>AA_AND2</type>
<position>78.5,-86.5</position>
<input>
<ID>IN_0</ID>807 </input>
<input>
<ID>IN_1</ID>809 </input>
<output>
<ID>OUT</ID>814 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>782</ID>
<type>DA_FROM</type>
<position>123.5,-111</position>
<input>
<ID>IN_0</ID>857 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B2</lparam></gate>
<gate>
<ID>757</ID>
<type>AE_OR2</type>
<position>85,-84.5</position>
<input>
<ID>IN_0</ID>812 </input>
<input>
<ID>IN_1</ID>814 </input>
<output>
<ID>OUT</ID>816 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>758</ID>
<type>DE_TO</type>
<position>117.5,-85</position>
<input>
<ID>IN_0</ID>591 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clrPC</lparam></gate>
<gate>
<ID>425</ID>
<type>AE_OR2</type>
<position>112.5,-85</position>
<input>
<ID>IN_0</ID>593 </input>
<input>
<ID>IN_1</ID>596 </input>
<output>
<ID>OUT</ID>591 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1118</ID>
<type>BE_JKFF_LOW</type>
<position>56,-20.5</position>
<input>
<ID>J</ID>1258 </input>
<input>
<ID>K</ID>1273 </input>
<output>
<ID>Q</ID>1243 </output>
<input>
<ID>clock</ID>1244 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>760</ID>
<type>DA_FROM</type>
<position>101.5,-83</position>
<input>
<ID>IN_0</ID>826 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>761</ID>
<type>DA_FROM</type>
<position>101.5,-85</position>
<input>
<ID>IN_0</ID>827 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T1</lparam></gate>
<gate>
<ID>287</ID>
<type>DM_NOR8</type>
<position>-43.5,-45.5</position>
<input>
<ID>IN_0</ID>383 </input>
<input>
<ID>IN_1</ID>385 </input>
<input>
<ID>IN_2</ID>381 </input>
<input>
<ID>IN_3</ID>386 </input>
<input>
<ID>IN_4</ID>388 </input>
<input>
<ID>IN_5</ID>382 </input>
<input>
<ID>IN_6</ID>387 </input>
<input>
<ID>IN_7</ID>384 </input>
<output>
<ID>OUT</ID>389 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>762</ID>
<type>AA_AND2</type>
<position>106.5,-84</position>
<input>
<ID>IN_0</ID>826 </input>
<input>
<ID>IN_1</ID>827 </input>
<output>
<ID>OUT</ID>593 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>763</ID>
<type>DE_TO</type>
<position>170.5,-102.5</position>
<input>
<ID>IN_0</ID>1020 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incPC</lparam></gate>
<gate>
<ID>1297</ID>
<type>DE_TO</type>
<position>-40.5,-144</position>
<input>
<ID>IN_0</ID>1369 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B8</lparam></gate>
<gate>
<ID>764</ID>
<type>DA_FROM</type>
<position>133.5,-81.5</position>
<input>
<ID>IN_0</ID>831 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>1117</ID>
<type>AE_OR2</type>
<position>40,-114</position>
<input>
<ID>IN_0</ID>1239 </input>
<input>
<ID>IN_1</ID>1240 </input>
<output>
<ID>OUT</ID>1242 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>784</ID>
<type>AE_SMALL_INVERTER</type>
<position>123.5,-113</position>
<input>
<ID>IN_0</ID>838 </input>
<output>
<ID>OUT_0</ID>1010 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>767</ID>
<type>DA_FROM</type>
<position>137.5,-83.5</position>
<input>
<ID>IN_0</ID>1023 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T1</lparam></gate>
<gate>
<ID>1101</ID>
<type>AA_LABEL</type>
<position>37.5,-98.5</position>
<gparam>LABEL_TEXT IEN Set/Reset</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>768</ID>
<type>DA_FROM</type>
<position>137.5,-87</position>
<input>
<ID>IN_0</ID>1024 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>769</ID>
<type>DA_FROM</type>
<position>137.5,-89</position>
<input>
<ID>IN_0</ID>1025 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T2</lparam></gate>
<gate>
<ID>770</ID>
<type>DA_FROM</type>
<position>137.5,-96.5</position>
<input>
<ID>IN_0</ID>1056 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>1106</ID>
<type>AA_AND2</type>
<position>40,-105.5</position>
<input>
<ID>IN_0</ID>1231 </input>
<input>
<ID>IN_1</ID>1232 </input>
<output>
<ID>OUT</ID>1230 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>771</ID>
<type>DA_FROM</type>
<position>137.5,-98.5</position>
<input>
<ID>IN_0</ID>1057 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T6</lparam></gate>
<gate>
<ID>772</ID>
<type>DA_FROM</type>
<position>119.5,-101</position>
<input>
<ID>IN_0</ID>833 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac15</lparam></gate>
<gate>
<ID>1080</ID>
<type>DA_FROM</type>
<position>18.5,-92</position>
<input>
<ID>IN_0</ID>1202 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID FGO</lparam></gate>
<gate>
<ID>773</ID>
<type>AE_SMALL_INVERTER</type>
<position>123.5,-101</position>
<input>
<ID>IN_0</ID>833 </input>
<output>
<ID>OUT_0</ID>848 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>775</ID>
<type>DA_FROM</type>
<position>123.5,-103</position>
<input>
<ID>IN_0</ID>850 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B4</lparam></gate>
<gate>
<ID>1109</ID>
<type>DA_FROM</type>
<position>35,-106.5</position>
<input>
<ID>IN_0</ID>1232 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B7</lparam></gate>
<gate>
<ID>776</ID>
<type>DA_FROM</type>
<position>123.5,-105</position>
<input>
<ID>IN_0</ID>851 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac15</lparam></gate>
<gate>
<ID>1114</ID>
<type>AA_AND2</type>
<position>32.5,-115.5</position>
<input>
<ID>IN_0</ID>1237 </input>
<input>
<ID>IN_1</ID>1238 </input>
<output>
<ID>OUT</ID>1240 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>779</ID>
<type>DA_FROM</type>
<position>123.5,-107</position>
<input>
<ID>IN_0</ID>853 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B3</lparam></gate>
<gate>
<ID>246</ID>
<type>FF_GND</type>
<position>258.5,-57.5</position>
<output>
<ID>OUT_0</ID>541 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>780</ID>
<type>DA_FROM</type>
<position>123.5,-109</position>
<input>
<ID>IN_0</ID>855 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC_zero</lparam></gate>
<gate>
<ID>781</ID>
<type>DA_FROM</type>
<position>123.5,-117</position>
<input>
<ID>IN_0</ID>1004 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>783</ID>
<type>DA_FROM</type>
<position>119.5,-113</position>
<input>
<ID>IN_0</ID>838 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID E</lparam></gate>
<gate>
<ID>1276</ID>
<type>DA_FROM</type>
<position>-44.5,-128</position>
<input>
<ID>IN_0</ID>1361 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir0</lparam></gate>
<gate>
<ID>785</ID>
<type>DA_FROM</type>
<position>123.5,-115</position>
<input>
<ID>IN_0</ID>1011 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B1</lparam></gate>
<gate>
<ID>788</ID>
<type>DA_FROM</type>
<position>125.5,-121.5</position>
<input>
<ID>IN_0</ID>1013 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID FGI</lparam></gate>
<gate>
<ID>790</ID>
<type>DA_FROM</type>
<position>125.5,-129.5</position>
<input>
<ID>IN_0</ID>1019 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>791</ID>
<type>DA_FROM</type>
<position>121.5,-125.5</position>
<input>
<ID>IN_0</ID>840 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID FGO</lparam></gate>
<gate>
<ID>1125</ID>
<type>AA_AND3</type>
<position>44,-17.5</position>
<input>
<ID>IN_0</ID>1271 </input>
<input>
<ID>IN_1</ID>1246 </input>
<input>
<ID>IN_2</ID>1247 </input>
<output>
<ID>OUT</ID>1258 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>792</ID>
<type>DA_FROM</type>
<position>125.5,-127.5</position>
<input>
<ID>IN_0</ID>1015 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B8</lparam></gate>
<gate>
<ID>1156</ID>
<type>AA_AND3</type>
<position>44,-23.5</position>
<input>
<ID>IN_0</ID>1247 </input>
<input>
<ID>IN_1</ID>1246 </input>
<input>
<ID>IN_2</ID>1272 </input>
<output>
<ID>OUT</ID>1273 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>793</ID>
<type>AE_SMALL_INVERTER</type>
<position>125.5,-125.5</position>
<input>
<ID>IN_0</ID>840 </input>
<output>
<ID>OUT_0</ID>1014 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>795</ID>
<type>AA_AND2</type>
<position>128.5,-102</position>
<input>
<ID>IN_0</ID>848 </input>
<input>
<ID>IN_1</ID>850 </input>
<output>
<ID>OUT</ID>1006 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>797</ID>
<type>AA_AND2</type>
<position>128.5,-106</position>
<input>
<ID>IN_0</ID>851 </input>
<input>
<ID>IN_1</ID>853 </input>
<output>
<ID>OUT</ID>1007 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>799</ID>
<type>AA_AND2</type>
<position>128.5,-110</position>
<input>
<ID>IN_0</ID>855 </input>
<input>
<ID>IN_1</ID>857 </input>
<output>
<ID>OUT</ID>1008 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1141</ID>
<type>BE_JKFF_LOW</type>
<position>22,-130</position>
<input>
<ID>J</ID>1261 </input>
<input>
<ID>K</ID>1262 </input>
<output>
<ID>Q</ID>1259 </output>
<input>
<ID>clock</ID>1260 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>808</ID>
<type>AE_OR4</type>
<position>135.5,-105</position>
<input>
<ID>IN_0</ID>1006 </input>
<input>
<ID>IN_1</ID>1007 </input>
<input>
<ID>IN_2</ID>1008 </input>
<input>
<ID>IN_3</ID>1009 </input>
<output>
<ID>OUT</ID>1005 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>812</ID>
<type>AA_AND2</type>
<position>130.5,-126.5</position>
<input>
<ID>IN_0</ID>1014 </input>
<input>
<ID>IN_1</ID>1015 </input>
<output>
<ID>OUT</ID>1030 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1149</ID>
<type>BE_JKFF_LOW</type>
<position>54,-130</position>
<input>
<ID>J</ID>1267 </input>
<input>
<ID>K</ID>1268 </input>
<output>
<ID>Q</ID>1265 </output>
<input>
<ID>clock</ID>1266 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>816</ID>
<type>AA_AND2</type>
<position>142.5,-124.5</position>
<input>
<ID>IN_0</ID>1029 </input>
<input>
<ID>IN_1</ID>1019 </input>
<output>
<ID>OUT</ID>1035 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>818</ID>
<type>DE_OR8</type>
<position>164.5,-102.5</position>
<input>
<ID>IN_0</ID>1031 </input>
<input>
<ID>IN_1</ID>1032 </input>
<input>
<ID>IN_2</ID>1058 </input>
<input>
<ID>IN_3</ID>1034 </input>
<input>
<ID>IN_4</ID>95 </input>
<input>
<ID>IN_5</ID>95 </input>
<input>
<ID>IN_6</ID>95 </input>
<input>
<ID>IN_7</ID>1035 </input>
<output>
<ID>OUT</ID>1020 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>820</ID>
<type>AA_AND2</type>
<position>142.5,-82.5</position>
<input>
<ID>IN_0</ID>1022 </input>
<input>
<ID>IN_1</ID>1023 </input>
<output>
<ID>OUT</ID>1031 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>822</ID>
<type>AA_AND2</type>
<position>142.5,-88</position>
<input>
<ID>IN_0</ID>1024 </input>
<input>
<ID>IN_1</ID>1025 </input>
<output>
<ID>OUT</ID>1032 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>826</ID>
<type>AE_OR2</type>
<position>136.5,-123.5</position>
<input>
<ID>IN_0</ID>1028 </input>
<input>
<ID>IN_1</ID>1030 </input>
<output>
<ID>OUT</ID>1029 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1034</ID>
<type>DA_FROM</type>
<position>16,-52</position>
<input>
<ID>IN_0</ID>1172 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac0</lparam></gate>
<gate>
<ID>827</ID>
<type>DE_TO</type>
<position>194,-85</position>
<input>
<ID>IN_0</ID>1043 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID busPC</lparam></gate>
<gate>
<ID>1165</ID>
<type>DA_FROM</type>
<position>-49,-22</position>
<input>
<ID>IN_0</ID>1291 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID I</lparam></gate>
<gate>
<ID>832</ID>
<type>DA_FROM</type>
<position>178,-84</position>
<input>
<ID>IN_0</ID>345 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T0</lparam></gate>
<gate>
<ID>833</ID>
<type>DA_FROM</type>
<position>178,-87.5</position>
<input>
<ID>IN_0</ID>1042 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>1139</ID>
<type>AA_LABEL</type>
<position>37,-122</position>
<gparam>LABEL_TEXT FGI/O Set/Reset</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>834</ID>
<type>DA_FROM</type>
<position>178,-89.5</position>
<input>
<ID>IN_0</ID>1041 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>1147</ID>
<type>DA_FROM</type>
<position>11,-132</position>
<input>
<ID>IN_0</ID>1263 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>1178</ID>
<type>AA_AND2</type>
<position>-36.5,-24</position>
<input>
<ID>IN_0</ID>1290 </input>
<input>
<ID>IN_1</ID>1287 </input>
<output>
<ID>OUT</ID>1289 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>843</ID>
<type>AA_AND2</type>
<position>183,-88.5</position>
<input>
<ID>IN_0</ID>1042 </input>
<input>
<ID>IN_1</ID>1041 </input>
<output>
<ID>OUT</ID>1045 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>846</ID>
<type>AA_LABEL</type>
<position>133,-137</position>
<gparam>LABEL_TEXT DR Commands</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>847</ID>
<type>AA_LABEL</type>
<position>37.5,-2.5</position>
<gparam>LABEL_TEXT Flip Flops</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1181</ID>
<type>AE_SMALL_INVERTER</type>
<position>-45,-23</position>
<input>
<ID>IN_0</ID>1291 </input>
<output>
<ID>OUT_0</ID>1290 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>848</ID>
<type>DE_TO</type>
<position>115.5,-149</position>
<input>
<ID>IN_0</ID>1050 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ldDR</lparam></gate>
<gate>
<ID>1</ID>
<type>AE_SMALL_INVERTER</type>
<position>88.5,-59</position>
<input>
<ID>IN_0</ID>148 </input>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1027</ID>
<type>DA_FROM</type>
<position>16,-36</position>
<input>
<ID>IN_0</ID>1167 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>850</ID>
<type>DA_FROM</type>
<position>98.5,-145</position>
<input>
<ID>IN_0</ID>1047 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>851</ID>
<type>DA_FROM</type>
<position>98.5,-147</position>
<input>
<ID>IN_0</ID>1048 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>852</ID>
<type>DA_FROM</type>
<position>98.5,-149</position>
<input>
<ID>IN_0</ID>1046 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>1032</ID>
<type>DA_FROM</type>
<position>16,-46</position>
<input>
<ID>IN_0</ID>1170 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac15</lparam></gate>
<gate>
<ID>853</ID>
<type>DA_FROM</type>
<position>98.5,-151</position>
<input>
<ID>IN_0</ID>1049 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>855</ID>
<type>AE_OR4</type>
<position>103.5,-148</position>
<input>
<ID>IN_0</ID>1047 </input>
<input>
<ID>IN_1</ID>1048 </input>
<input>
<ID>IN_2</ID>1046 </input>
<input>
<ID>IN_3</ID>1049 </input>
<output>
<ID>OUT</ID>1052 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>857</ID>
<type>AA_AND2</type>
<position>110.5,-149</position>
<input>
<ID>IN_0</ID>1052 </input>
<input>
<ID>IN_1</ID>1051 </input>
<output>
<ID>OUT</ID>1050 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1035</ID>
<type>DA_FROM</type>
<position>16,-48</position>
<input>
<ID>IN_0</ID>1174 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>858</ID>
<type>DA_FROM</type>
<position>98.5,-153</position>
<input>
<ID>IN_0</ID>1051 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>1194</ID>
<type>DA_FROM</type>
<position>-48.5,-34</position>
<input>
<ID>IN_0</ID>357 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr0</lparam></gate>
<gate>
<ID>859</ID>
<type>DE_TO</type>
<position>136.5,-149</position>
<input>
<ID>IN_0</ID>1055 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incDR</lparam></gate>
<gate>
<ID>860</ID>
<type>DA_FROM</type>
<position>126.5,-148</position>
<input>
<ID>IN_0</ID>1053 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>1040</ID>
<type>AA_AND3</type>
<position>21,-44</position>
<input>
<ID>IN_0</ID>1171 </input>
<input>
<ID>IN_1</ID>1169 </input>
<input>
<ID>IN_2</ID>1170 </input>
<output>
<ID>OUT</ID>1177 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>861</ID>
<type>DA_FROM</type>
<position>126.5,-150</position>
<input>
<ID>IN_0</ID>1054 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>862</ID>
<type>AA_AND2</type>
<position>131.5,-149</position>
<input>
<ID>IN_0</ID>1053 </input>
<input>
<ID>IN_1</ID>1054 </input>
<output>
<ID>OUT</ID>1055 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1197</ID>
<type>DA_FROM</type>
<position>-56,-37</position>
<input>
<ID>IN_0</ID>361 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr3</lparam></gate>
<gate>
<ID>864</ID>
<type>AA_AND3</type>
<position>142.5,-96.5</position>
<input>
<ID>IN_0</ID>1059 </input>
<input>
<ID>IN_1</ID>1056 </input>
<input>
<ID>IN_2</ID>1057 </input>
<output>
<ID>OUT</ID>1058 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>1228</ID>
<type>DA_FROM</type>
<position>-56,-56.5</position>
<input>
<ID>IN_0</ID>428 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac5</lparam></gate>
<gate>
<ID>865</ID>
<type>DA_FROM</type>
<position>137.5,-94.5</position>
<input>
<ID>IN_0</ID>1059 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR_zero</lparam></gate>
<gate>
<ID>1043</ID>
<type>AE_OR3</type>
<position>36,-44</position>
<input>
<ID>IN_0</ID>1176 </input>
<input>
<ID>IN_1</ID>1177 </input>
<input>
<ID>IN_2</ID>1178 </input>
<output>
<ID>OUT</ID>1185 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>866</ID>
<type>DE_TO</type>
<position>171,-149</position>
<input>
<ID>IN_0</ID>1060 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID busDR</lparam></gate>
<gate>
<ID>1202</ID>
<type>DA_FROM</type>
<position>-48.5,-42</position>
<input>
<ID>IN_0</ID>383 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr8</lparam></gate>
<gate>
<ID>867</ID>
<type>DA_FROM</type>
<position>155,-151</position>
<input>
<ID>IN_0</ID>1064 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>868</ID>
<type>DA_FROM</type>
<position>155,-153</position>
<input>
<ID>IN_0</ID>1065 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T6</lparam></gate>
<gate>
<ID>869</ID>
<type>DA_FROM</type>
<position>153,-145</position>
<input>
<ID>IN_0</ID>1062 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>870</ID>
<type>DA_FROM</type>
<position>153,-147</position>
<input>
<ID>IN_0</ID>1063 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>1205</ID>
<type>DA_FROM</type>
<position>-56,-45</position>
<input>
<ID>IN_0</ID>386 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr11</lparam></gate>
<gate>
<ID>872</ID>
<type>AE_OR2</type>
<position>166,-149</position>
<input>
<ID>IN_0</ID>1069 </input>
<input>
<ID>IN_1</ID>1068 </input>
<output>
<ID>OUT</ID>1060 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>874</ID>
<type>AA_AND2</type>
<position>160,-146</position>
<input>
<ID>IN_0</ID>1062 </input>
<input>
<ID>IN_1</ID>1063 </input>
<output>
<ID>OUT</ID>1069 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1210</ID>
<type>DA_FROM</type>
<position>-48.5,-51.5</position>
<input>
<ID>IN_0</ID>391 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac0</lparam></gate>
<gate>
<ID>875</ID>
<type>AA_AND2</type>
<position>160,-152</position>
<input>
<ID>IN_0</ID>1064 </input>
<input>
<ID>IN_1</ID>1065 </input>
<output>
<ID>OUT</ID>1068 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>876</ID>
<type>AA_LABEL</type>
<position>134,-163.5</position>
<gparam>LABEL_TEXT IR Commands</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1056</ID>
<type>AA_AND2</type>
<position>46,-49.5</position>
<input>
<ID>IN_0</ID>1191 </input>
<input>
<ID>IN_1</ID>351 </input>
<output>
<ID>OUT</ID>1194 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>877</ID>
<type>DE_TO</type>
<position>123.5,-173</position>
<input>
<ID>IN_0</ID>1073 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ldIR</lparam></gate>
<gate>
<ID>878</ID>
<type>DA_FROM</type>
<position>109.5,-172</position>
<input>
<ID>IN_0</ID>1070 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>879</ID>
<type>AE_SMALL_INVERTER</type>
<position>113.5,-172</position>
<input>
<ID>IN_0</ID>1070 </input>
<output>
<ID>OUT_0</ID>1072 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>880</ID>
<type>DA_FROM</type>
<position>113.5,-174</position>
<input>
<ID>IN_0</ID>1071 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T1</lparam></gate>
<gate>
<ID>1244</ID>
<type>DE_TO</type>
<position>-38,-95</position>
<input>
<ID>IN_0</ID>1349 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INPR</lparam></gate>
<gate>
<ID>881</ID>
<type>AA_AND2</type>
<position>118.5,-173</position>
<input>
<ID>IN_0</ID>1072 </input>
<input>
<ID>IN_1</ID>1071 </input>
<output>
<ID>OUT</ID>1073 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1059</ID>
<type>AA_LABEL</type>
<position>38,-76.5</position>
<gparam>LABEL_TEXT R Set/Reset</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>882</ID>
<type>DA_FROM</type>
<position>139.5,-172</position>
<input>
<ID>IN_0</ID>1074 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>884</ID>
<type>DA_FROM</type>
<position>143.5,-174</position>
<input>
<ID>IN_0</ID>1075 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T2</lparam></gate>
<gate>
<ID>1064</ID>
<type>DA_FROM</type>
<position>20.5,-81.5</position>
<input>
<ID>IN_0</ID>1198 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T0</lparam></gate>
<gate>
<ID>885</ID>
<type>AA_AND2</type>
<position>148.5,-173</position>
<input>
<ID>IN_0</ID>1076 </input>
<input>
<ID>IN_1</ID>1075 </input>
<output>
<ID>OUT</ID>1077 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>886</ID>
<type>DE_TO</type>
<position>153.5,-173</position>
<input>
<ID>IN_0</ID>1077 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID busIR</lparam></gate>
<gate>
<ID>1093</ID>
<type>DA_FROM</type>
<position>16,-63</position>
<input>
<ID>IN_0</ID>1211 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>888</ID>
<type>AA_LABEL</type>
<position>134,-183</position>
<gparam>LABEL_TEXT TR Commands</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>889</ID>
<type>DE_TO</type>
<position>123.5,-193</position>
<input>
<ID>IN_0</ID>1081 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ldTR</lparam></gate>
<gate>
<ID>890</ID>
<type>DA_FROM</type>
<position>113.5,-192</position>
<input>
<ID>IN_0</ID>1086 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>892</ID>
<type>DA_FROM</type>
<position>113.5,-194</position>
<input>
<ID>IN_0</ID>1079 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T0</lparam></gate>
<gate>
<ID>1072</ID>
<type>DA_FROM</type>
<position>24.5,-87.5</position>
<input>
<ID>IN_0</ID>1222 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IEN</lparam></gate>
<gate>
<ID>893</ID>
<type>AA_AND2</type>
<position>118.5,-193</position>
<input>
<ID>IN_0</ID>1086 </input>
<input>
<ID>IN_1</ID>1079 </input>
<output>
<ID>OUT</ID>1081 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>894</ID>
<type>DA_FROM</type>
<position>143.5,-192</position>
<input>
<ID>IN_0</ID>1087 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>895</ID>
<type>DA_FROM</type>
<position>143.5,-194</position>
<input>
<ID>IN_0</ID>1083 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T1</lparam></gate>
<gate>
<ID>1229</ID>
<type>DA_FROM</type>
<position>-48.5,-57.5</position>
<input>
<ID>IN_0</ID>390 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac6</lparam></gate>
<gate>
<ID>896</ID>
<type>AA_AND2</type>
<position>148.5,-193</position>
<input>
<ID>IN_0</ID>1087 </input>
<input>
<ID>IN_1</ID>1083 </input>
<output>
<ID>OUT</ID>1085 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>897</ID>
<type>DE_TO</type>
<position>153.5,-193</position>
<input>
<ID>IN_0</ID>1085 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID busTR</lparam></gate>
<gate>
<ID>39</ID>
<type>AA_AND2</type>
<position>21,-68</position>
<input>
<ID>IN_0</ID>349 </input>
<input>
<ID>IN_1</ID>350 </input>
<output>
<ID>OUT</ID>355 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1203</ID>
<type>DA_FROM</type>
<position>-56,-43</position>
<input>
<ID>IN_0</ID>385 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr9</lparam></gate>
<gate>
<ID>898</ID>
<type>AA_LABEL</type>
<position>134,-202.5</position>
<gparam>LABEL_TEXT AC Commands</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1208</ID>
<type>DA_FROM</type>
<position>-48.5,-48</position>
<input>
<ID>IN_0</ID>382 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr14</lparam></gate>
<gate>
<ID>901</ID>
<type>DA_FROM</type>
<position>82,-202</position>
<input>
<ID>IN_0</ID>1088 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>902</ID>
<type>DA_FROM</type>
<position>82,-204</position>
<input>
<ID>IN_0</ID>1089 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>1237</ID>
<type>DA_FROM</type>
<position>-48.5,-65.5</position>
<input>
<ID>IN_0</ID>562 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac14</lparam></gate>
<gate>
<ID>904</ID>
<type>DA_FROM</type>
<position>82,-208.5</position>
<input>
<ID>IN_0</ID>1092 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>905</ID>
<type>DA_FROM</type>
<position>82,-206</position>
<input>
<ID>IN_0</ID>1090 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>1242</ID>
<type>DE_TO</type>
<position>-38,-86</position>
<input>
<ID>IN_0</ID>1345 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>907</ID>
<type>DA_FROM</type>
<position>82,-218</position>
<input>
<ID>IN_0</ID>1097 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>1057</ID>
<type>DA_FROM</type>
<position>48,-46</position>
<input>
<ID>IN_0</ID>1195 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>908</ID>
<type>DA_FROM</type>
<position>82,-215.5</position>
<input>
<ID>IN_0</ID>1095 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B9</lparam></gate>
<gate>
<ID>910</ID>
<type>DA_FROM</type>
<position>82,-213.5</position>
<input>
<ID>IN_0</ID>1094 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B7</lparam></gate>
<gate>
<ID>1245</ID>
<type>DE_TO</type>
<position>-38,-101.5</position>
<input>
<ID>IN_0</ID>1352 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID COM</lparam></gate>
<gate>
<ID>912</ID>
<type>DA_FROM</type>
<position>82,-211.5</position>
<input>
<ID>IN_0</ID>1093 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B6</lparam></gate>
<gate>
<ID>913</ID>
<type>DA_FROM</type>
<position>88,-221.5</position>
<input>
<ID>IN_0</ID>1099 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>1091</ID>
<type>DA_FROM</type>
<position>16,-61</position>
<input>
<ID>IN_0</ID>1209 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B6</lparam></gate>
<gate>
<ID>914</ID>
<type>DA_FROM</type>
<position>88,-223.5</position>
<input>
<ID>IN_0</ID>1098 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B11</lparam></gate>
<gate>
<ID>1065</ID>
<type>DA_FROM</type>
<position>20.5,-83.5</position>
<input>
<ID>IN_0</ID>1199 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T1</lparam></gate>
<gate>
<ID>916</ID>
<type>AE_OR3</type>
<position>87,-204</position>
<input>
<ID>IN_0</ID>1088 </input>
<input>
<ID>IN_1</ID>1089 </input>
<input>
<ID>IN_2</ID>1090 </input>
<output>
<ID>OUT</ID>1091 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>918</ID>
<type>AA_AND2</type>
<position>93,-205.5</position>
<input>
<ID>IN_0</ID>1091 </input>
<input>
<ID>IN_1</ID>1092 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1253</ID>
<type>AA_AND2</type>
<position>-43,-86</position>
<input>
<ID>IN_0</ID>1343 </input>
<input>
<ID>IN_1</ID>1344 </input>
<output>
<ID>OUT</ID>1345 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>920</ID>
<type>AE_OR3</type>
<position>87,-213.5</position>
<input>
<ID>IN_0</ID>1093 </input>
<input>
<ID>IN_1</ID>1094 </input>
<input>
<ID>IN_2</ID>1095 </input>
<output>
<ID>OUT</ID>1096 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>922</ID>
<type>AA_AND2</type>
<position>93,-214.5</position>
<input>
<ID>IN_0</ID>1096 </input>
<input>
<ID>IN_1</ID>1097 </input>
<output>
<ID>OUT</ID>1100 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>924</ID>
<type>AA_AND2</type>
<position>93,-222.5</position>
<input>
<ID>IN_0</ID>1099 </input>
<input>
<ID>IN_1</ID>1098 </input>
<output>
<ID>OUT</ID>1102 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>926</ID>
<type>AE_OR3</type>
<position>99,-214.5</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>1100 </input>
<input>
<ID>IN_2</ID>1102 </input>
<output>
<ID>OUT</ID>1103 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>927</ID>
<type>DE_TO</type>
<position>134,-215</position>
<input>
<ID>IN_0</ID>153 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clrAC</lparam></gate>
<gate>
<ID>929</ID>
<type>AA_AND2</type>
<position>123,-214</position>
<input>
<ID>IN_0</ID>1105 </input>
<input>
<ID>IN_1</ID>1106 </input>
<output>
<ID>OUT</ID>333 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>930</ID>
<type>DA_FROM</type>
<position>118,-213</position>
<input>
<ID>IN_0</ID>1105 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>1266</ID>
<type>DA_FROM</type>
<position>-54,-103.5</position>
<input>
<ID>IN_0</ID>1354 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>931</ID>
<type>DA_FROM</type>
<position>118,-215</position>
<input>
<ID>IN_0</ID>1106 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B11</lparam></gate>
<gate>
<ID>932</ID>
<type>DE_TO</type>
<position>157.5,-215</position>
<input>
<ID>IN_0</ID>1109 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID incAC</lparam></gate>
<gate>
<ID>1294</ID>
<type>DE_TO</type>
<position>-40.5,-138</position>
<input>
<ID>IN_0</ID>1366 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B5</lparam></gate>
<gate>
<ID>1269</ID>
<type>AA_AND2</type>
<position>-43,-108</position>
<input>
<ID>IN_0</ID>1356 </input>
<input>
<ID>IN_1</ID>1357 </input>
<output>
<ID>OUT</ID>1355 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>936</ID>
<type>DA_FROM</type>
<position>147.5,-214</position>
<input>
<ID>IN_0</ID>1107 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>937</ID>
<type>DA_FROM</type>
<position>147.5,-216</position>
<input>
<ID>IN_0</ID>1108 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B5</lparam></gate>
<gate>
<ID>1115</ID>
<type>DA_FROM</type>
<position>27.5,-116.5</position>
<input>
<ID>IN_0</ID>1238 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T2</lparam></gate>
<gate>
<ID>938</ID>
<type>DE_TO</type>
<position>189.5,-215</position>
<input>
<ID>IN_0</ID>1110 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID busAC</lparam></gate>
<gate>
<ID>940</ID>
<type>AE_OR2</type>
<position>184.5,-215</position>
<input>
<ID>IN_0</ID>1116 </input>
<input>
<ID>IN_1</ID>1113 </input>
<output>
<ID>OUT</ID>1110 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1120</ID>
<type>DA_FROM</type>
<position>28,-20.5</position>
<input>
<ID>IN_0</ID>1245 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>941</ID>
<type>DA_FROM</type>
<position>173.5,-216</position>
<input>
<ID>IN_0</ID>1112 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>942</ID>
<type>DA_FROM</type>
<position>173.5,-218</position>
<input>
<ID>IN_0</ID>1111 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B10</lparam></gate>
<gate>
<ID>1293</ID>
<type>DE_TO</type>
<position>-40.5,-136</position>
<input>
<ID>IN_0</ID>1365 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B4</lparam></gate>
<gate>
<ID>943</ID>
<type>AA_AND2</type>
<position>178.5,-217</position>
<input>
<ID>IN_0</ID>1112 </input>
<input>
<ID>IN_1</ID>1111 </input>
<output>
<ID>OUT</ID>1113 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1123</ID>
<type>AE_SMALL_INVERTER</type>
<position>32,-20.5</position>
<input>
<ID>IN_0</ID>1245 </input>
<output>
<ID>OUT_0</ID>1246 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>946</ID>
<type>DA_FROM</type>
<position>173.5,-212</position>
<input>
<ID>IN_0</ID>1115 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>1154</ID>
<type>AA_AND2</type>
<position>48,-133</position>
<input>
<ID>IN_0</ID>1269 </input>
<input>
<ID>IN_1</ID>1270 </input>
<output>
<ID>OUT</ID>1268 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>947</ID>
<type>DA_FROM</type>
<position>173.5,-214</position>
<input>
<ID>IN_0</ID>1114 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>948</ID>
<type>AA_AND2</type>
<position>178.5,-213</position>
<input>
<ID>IN_0</ID>1115 </input>
<input>
<ID>IN_1</ID>1114 </input>
<output>
<ID>OUT</ID>1116 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>950</ID>
<type>AA_LABEL</type>
<position>-109,-35</position>
<gparam>LABEL_TEXT ldOUTR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>951</ID>
<type>DE_TO</type>
<position>-106.5,-41</position>
<input>
<ID>IN_0</ID>1119 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ldOUTR</lparam></gate>
<gate>
<ID>952</ID>
<type>DA_FROM</type>
<position>-116.5,-40</position>
<input>
<ID>IN_0</ID>1118 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>953</ID>
<type>DA_FROM</type>
<position>-116.5,-42</position>
<input>
<ID>IN_0</ID>1117 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B10</lparam></gate>
<gate>
<ID>954</ID>
<type>AA_AND2</type>
<position>-111.5,-41</position>
<input>
<ID>IN_0</ID>1118 </input>
<input>
<ID>IN_1</ID>1117 </input>
<output>
<ID>OUT</ID>1119 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>955</ID>
<type>EE_VDD</type>
<position>219,-19.5</position>
<output>
<ID>OUT_0</ID>600 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>958</ID>
<type>DA_FROM</type>
<position>219.5,-31.5</position>
<input>
<ID>IN_0</ID>1136 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID clrSC</lparam></gate>
<gate>
<ID>959</ID>
<type>DE_TO</type>
<position>230.5,-24.5</position>
<input>
<ID>IN_0</ID>1129 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T2</lparam></gate>
<gate>
<ID>1291</ID>
<type>DE_TO</type>
<position>-40.5,-132</position>
<input>
<ID>IN_0</ID>1363 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B2</lparam></gate>
<gate>
<ID>961</ID>
<type>DE_TO</type>
<position>230.5,-26.5</position>
<input>
<ID>IN_0</ID>1127 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T0</lparam></gate>
<gate>
<ID>1300</ID>
<type>DE_TO</type>
<position>-40.5,-150</position>
<input>
<ID>IN_0</ID>1372 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B11</lparam></gate>
<gate>
<ID>1267</ID>
<type>DA_FROM</type>
<position>-48,-107</position>
<input>
<ID>IN_0</ID>1356 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>962</ID>
<type>DE_TO</type>
<position>235.5,-25.5</position>
<input>
<ID>IN_0</ID>1128 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T1</lparam></gate>
<gate>
<ID>963</ID>
<type>DE_TO</type>
<position>235.5,-23.5</position>
<input>
<ID>IN_0</ID>1130 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T3</lparam></gate>
<gate>
<ID>1272</ID>
<type>DA_FROM</type>
<position>-48,-113</position>
<input>
<ID>IN_0</ID>1358 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>965</ID>
<type>DE_TO</type>
<position>235.5,-21.5</position>
<input>
<ID>IN_0</ID>1132 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>966</ID>
<type>DE_TO</type>
<position>230.5,-20.5</position>
<input>
<ID>IN_0</ID>1133 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T6</lparam></gate>
<gate>
<ID>1086</ID>
<type>AA_AND2</type>
<position>21,-64</position>
<input>
<ID>IN_0</ID>1211 </input>
<input>
<ID>IN_1</ID>1212 </input>
<output>
<ID>OUT</ID>354 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>967</ID>
<type>DE_TO</type>
<position>235.5,-19.5</position>
<input>
<ID>IN_0</ID>1134 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T7</lparam></gate>
<gate>
<ID>1299</ID>
<type>DE_TO</type>
<position>-40.5,-148</position>
<input>
<ID>IN_0</ID>1371 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B10</lparam></gate>
<gate>
<ID>969</ID>
<type>BE_DECODER_3x8</type>
<position>225.5,-23</position>
<input>
<ID>ENABLE</ID>1135 </input>
<input>
<ID>IN_0</ID>1125 </input>
<input>
<ID>IN_1</ID>1126 </input>
<input>
<ID>IN_2</ID>1124 </input>
<output>
<ID>OUT_0</ID>1127 </output>
<output>
<ID>OUT_1</ID>1128 </output>
<output>
<ID>OUT_2</ID>1129 </output>
<output>
<ID>OUT_3</ID>1130 </output>
<output>
<ID>OUT_4</ID>1131 </output>
<output>
<ID>OUT_5</ID>1132 </output>
<output>
<ID>OUT_6</ID>1133 </output>
<output>
<ID>OUT_7</ID>1134 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>970</ID>
<type>AA_LABEL</type>
<position>223.5,-13</position>
<gparam>LABEL_TEXT Counter</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1121</ID>
<type>DA_FROM</type>
<position>39,-20.5</position>
<input>
<ID>IN_0</ID>1247 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T2</lparam></gate>
<gate>
<ID>972</ID>
<type>AA_LABEL</type>
<position>253,-3.5</position>
<gparam>LABEL_TEXT SC Commands</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1152</ID>
<type>DE_TO</type>
<position>59,-128</position>
<input>
<ID>IN_0</ID>1265 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID FGO</lparam></gate>
<gate>
<ID>973</ID>
<type>DE_TO</type>
<position>267.5,-52</position>
<input>
<ID>IN_0</ID>1152 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clrSC</lparam></gate>
<gate>
<ID>975</ID>
<type>DA_FROM</type>
<position>235.5,-41</position>
<input>
<ID>IN_0</ID>1149 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>977</ID>
<type>DA_FROM</type>
<position>235.5,-43</position>
<input>
<ID>IN_0</ID>1148 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T2</lparam></gate>
<gate>
<ID>1155</ID>
<type>DA_FROM</type>
<position>43,-134</position>
<input>
<ID>IN_0</ID>1270 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B10</lparam></gate>
<gate>
<ID>978</ID>
<type>DA_FROM</type>
<position>228.5,-45.5</position>
<input>
<ID>IN_0</ID>1138 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>982</ID>
<type>DA_FROM</type>
<position>228.5,-47.5</position>
<input>
<ID>IN_0</ID>1139 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>984</ID>
<type>DA_FROM</type>
<position>228.5,-49.5</position>
<input>
<ID>IN_0</ID>1137 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>986</ID>
<type>DA_FROM</type>
<position>229.5,-56</position>
<input>
<ID>IN_0</ID>1144 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>988</ID>
<type>DA_FROM</type>
<position>229.5,-58</position>
<input>
<ID>IN_0</ID>1145 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>989</ID>
<type>DA_FROM</type>
<position>229.5,-60</position>
<input>
<ID>IN_0</ID>1147 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>990</ID>
<type>DA_FROM</type>
<position>228.5,-53.5</position>
<input>
<ID>IN_0</ID>1143 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>298</ID>
<type>BB_CLOCK</type>
<position>260.5,-35.5</position>
<output>
<ID>CLK</ID>565 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 20</lparam></gate>
<gate>
<ID>992</ID>
<type>DA_FROM</type>
<position>235.5,-62.5</position>
<input>
<ID>IN_0</ID>1150 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>993</ID>
<type>DA_FROM</type>
<position>235.5,-64.5</position>
<input>
<ID>IN_0</ID>1151 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T6</lparam></gate>
<gate>
<ID>994</ID>
<type>DA_FROM</type>
<position>241.5,-67</position>
<input>
<ID>IN_0</ID>1157 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>1176</ID>
<type>AA_AND2</type>
<position>-36.5,-20</position>
<input>
<ID>IN_0</ID>1287 </input>
<input>
<ID>IN_1</ID>1291 </input>
<output>
<ID>OUT</ID>1284 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>997</ID>
<type>AE_OR4</type>
<position>233.5,-48.5</position>
<input>
<ID>IN_0</ID>1138 </input>
<input>
<ID>IN_1</ID>1139 </input>
<input>
<ID>IN_2</ID>1137 </input>
<input>
<ID>IN_3</ID>1140 </input>
<output>
<ID>OUT</ID>1141 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>999</ID>
<type>AA_AND2</type>
<position>240.5,-49.5</position>
<input>
<ID>IN_0</ID>1141 </input>
<input>
<ID>IN_1</ID>1143 </input>
<output>
<ID>OUT</ID>1154 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1007</ID>
<type>AA_AND2</type>
<position>240.5,-42</position>
<input>
<ID>IN_0</ID>1149 </input>
<input>
<ID>IN_1</ID>1148 </input>
<output>
<ID>OUT</ID>1153 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1009</ID>
<type>AA_AND2</type>
<position>240.5,-63.5</position>
<input>
<ID>IN_0</ID>1150 </input>
<input>
<ID>IN_1</ID>1151 </input>
<output>
<ID>OUT</ID>1156 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1011</ID>
<type>DE_OR8</type>
<position>261.5,-52</position>
<input>
<ID>IN_0</ID>1153 </input>
<input>
<ID>IN_1</ID>1154 </input>
<input>
<ID>IN_2</ID>1155 </input>
<input>
<ID>IN_3</ID>1156 </input>
<input>
<ID>IN_4</ID>541 </input>
<input>
<ID>IN_5</ID>587 </input>
<input>
<ID>IN_6</ID>1158 </input>
<input>
<ID>IN_7</ID>1157 </input>
<output>
<ID>OUT</ID>1152 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1033</ID>
<type>DA_FROM</type>
<position>16,-50</position>
<input>
<ID>IN_0</ID>1173 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B7</lparam></gate>
<gate>
<ID>1012</ID>
<type>AA_LABEL</type>
<position>265,-12</position>
<gparam>LABEL_TEXT START/HALT Command</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1013</ID>
<type>DE_TO</type>
<position>272.5,-21.5</position>
<input>
<ID>IN_0</ID>96 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID S</lparam></gate>
<gate>
<ID>1016</ID>
<type>DA_FROM</type>
<position>244.5,-23.5</position>
<input>
<ID>IN_0</ID>151 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>1041</ID>
<type>AA_AND3</type>
<position>21,-50</position>
<input>
<ID>IN_0</ID>1174 </input>
<input>
<ID>IN_1</ID>1173 </input>
<input>
<ID>IN_2</ID>1172 </input>
<output>
<ID>OUT</ID>1178 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>1020</ID>
<type>DA_FROM</type>
<position>22,-20.5</position>
<input>
<ID>IN_0</ID>1271 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir15</lparam></gate>
<gate>
<ID>310</ID>
<type>DE_TO</type>
<position>277,-36.5</position>
<input>
<ID>IN_0</ID>563 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>1025</ID>
<type>DE_TO</type>
<position>58,-44</position>
<input>
<ID>IN_0</ID>1165 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID E</lparam></gate>
<gate>
<ID>1029</ID>
<type>DA_FROM</type>
<position>16,-40</position>
<input>
<ID>IN_0</ID>1168 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Cout</lparam></gate>
<gate>
<ID>1031</ID>
<type>DA_FROM</type>
<position>16,-42</position>
<input>
<ID>IN_0</ID>1171 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>147</ID>
<type>DA_FROM</type>
<position>124,-218.5</position>
<input>
<ID>IN_0</ID>344 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID START</lparam></gate>
<gate>
<ID>1037</ID>
<type>BE_JKFF_LOW</type>
<position>53,-46</position>
<input>
<ID>J</ID>1185 </input>
<input>
<ID>K</ID>1194 </input>
<output>
<ID>Q</ID>1165 </output>
<input>
<ID>clock</ID>1195 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1039</ID>
<type>AA_AND3</type>
<position>21,-38</position>
<input>
<ID>IN_0</ID>1167 </input>
<input>
<ID>IN_1</ID>1166 </input>
<input>
<ID>IN_2</ID>1168 </input>
<output>
<ID>OUT</ID>1176 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>367</ID>
<type>AA_LABEL</type>
<position>249,-30.5</position>
<gparam>LABEL_TEXT MANUAL HALT</gparam>
<gparam>TEXT_HEIGHT 0.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1052</ID>
<type>AE_SMALL_INVERTER</type>
<position>41,-48.5</position>
<input>
<ID>IN_0</ID>1185 </input>
<output>
<ID>OUT_0</ID>1191 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1058</ID>
<type>BE_JKFF_LOW</type>
<position>49.5,-87</position>
<input>
<ID>J</ID>1213 </input>
<input>
<ID>K</ID>1227 </input>
<output>
<ID>Q</ID>1196 </output>
<input>
<ID>clock</ID>1197 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>375</ID>
<type>DA_FROM</type>
<position>241.5,-71</position>
<input>
<ID>IN_0</ID>587 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID START</lparam></gate>
<gate>
<ID>1060</ID>
<type>DE_TO</type>
<position>54.5,-85</position>
<input>
<ID>IN_0</ID>1196 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>1066</ID>
<type>DA_FROM</type>
<position>20.5,-85.5</position>
<input>
<ID>IN_0</ID>1200 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T2</lparam></gate>
<gate>
<ID>1068</ID>
<type>AE_SMALL_INVERTER</type>
<position>24.5,-81.5</position>
<input>
<ID>IN_0</ID>1198 </input>
<output>
<ID>OUT_0</ID>1219 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1076</ID>
<type>AE_OR2</type>
<position>23.5,-91</position>
<input>
<ID>IN_0</ID>1201 </input>
<input>
<ID>IN_1</ID>1202 </input>
<output>
<ID>OUT</ID>1223 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1078</ID>
<type>DA_FROM</type>
<position>18.5,-90</position>
<input>
<ID>IN_0</ID>1201 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID FGI</lparam></gate>
<gate>
<ID>1082</ID>
<type>AA_AND2</type>
<position>21,-56</position>
<input>
<ID>IN_0</ID>1208 </input>
<input>
<ID>IN_1</ID>1207 </input>
<output>
<ID>OUT</ID>352 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1084</ID>
<type>AA_AND2</type>
<position>21,-60</position>
<input>
<ID>IN_0</ID>1210 </input>
<input>
<ID>IN_1</ID>1209 </input>
<output>
<ID>OUT</ID>353 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1087</ID>
<type>DA_FROM</type>
<position>16,-57</position>
<input>
<ID>IN_0</ID>1207 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>1088</ID>
<type>DA_FROM</type>
<position>16,-55</position>
<input>
<ID>IN_0</ID>1208 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>1092</ID>
<type>DA_FROM</type>
<position>16,-59</position>
<input>
<ID>IN_0</ID>1210 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>1094</ID>
<type>DA_FROM</type>
<position>16,-65</position>
<input>
<ID>IN_0</ID>1212 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B7</lparam></gate>
<gate>
<ID>1096</ID>
<type>DA_AND8</type>
<position>32,-85</position>
<input>
<ID>IN_0</ID>1219 </input>
<input>
<ID>IN_1</ID>1220 </input>
<input>
<ID>IN_2</ID>1221 </input>
<input>
<ID>IN_3</ID>1222 </input>
<input>
<ID>IN_4</ID>1223 </input>
<output>
<ID>OUT</ID>1213 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1097</ID>
<type>DA_FROM</type>
<position>38.5,-93</position>
<input>
<ID>IN_0</ID>1224 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T2</lparam></gate>
<gate>
<ID>1098</ID>
<type>DA_FROM</type>
<position>38.5,-91</position>
<input>
<ID>IN_0</ID>1225 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>1102</ID>
<type>DA_FROM</type>
<position>41,-110</position>
<input>
<ID>IN_0</ID>1229 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>1103</ID>
<type>BE_JKFF_LOW</type>
<position>46,-110</position>
<input>
<ID>J</ID>1230 </input>
<input>
<ID>K</ID>1242 </input>
<output>
<ID>Q</ID>1228 </output>
<input>
<ID>clock</ID>1229 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1104</ID>
<type>DE_TO</type>
<position>51,-108</position>
<input>
<ID>IN_0</ID>1228 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IEN</lparam></gate>
<gate>
<ID>1108</ID>
<type>DA_FROM</type>
<position>35,-104.5</position>
<input>
<ID>IN_0</ID>1231 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>1111</ID>
<type>DA_FROM</type>
<position>27.5,-110.5</position>
<input>
<ID>IN_0</ID>1233 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>1119</ID>
<type>DA_FROM</type>
<position>51,-20.5</position>
<input>
<ID>IN_0</ID>1244 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>1138</ID>
<type>AA_LABEL</type>
<position>37.5,-10</position>
<gparam>LABEL_TEXT I Set/Reset</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1140</ID>
<type>DA_FROM</type>
<position>17,-130</position>
<input>
<ID>IN_0</ID>1260 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>1142</ID>
<type>DE_TO</type>
<position>27,-128</position>
<input>
<ID>IN_0</ID>1259 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID FGI</lparam></gate>
<gate>
<ID>1144</ID>
<type>AA_TOGGLE</type>
<position>17,-128</position>
<output>
<ID>OUT_0</ID>1261 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1146</ID>
<type>AA_AND2</type>
<position>16,-133</position>
<input>
<ID>IN_0</ID>1263 </input>
<input>
<ID>IN_1</ID>1264 </input>
<output>
<ID>OUT</ID>1262 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>335</ID>
<type>AE_OR2</type>
<position>266,-40</position>
<input>
<ID>IN_0</ID>569 </input>
<input>
<ID>IN_1</ID>572 </input>
<output>
<ID>OUT</ID>574 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1148</ID>
<type>DA_FROM</type>
<position>11,-134</position>
<input>
<ID>IN_0</ID>1264 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B11</lparam></gate>
<gate>
<ID>1150</ID>
<type>DA_FROM</type>
<position>43,-132</position>
<input>
<ID>IN_0</ID>1269 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>1153</ID>
<type>AA_TOGGLE</type>
<position>49,-128</position>
<output>
<ID>OUT_0</ID>1267 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1158</ID>
<type>AE_SMALL_INVERTER</type>
<position>26,-25.5</position>
<input>
<ID>IN_0</ID>1271 </input>
<output>
<ID>OUT_0</ID>1272 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1159</ID>
<type>AA_LABEL</type>
<position>-105.5,-1.5</position>
<gparam>LABEL_TEXT Misc.</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>1160</ID>
<type>AA_LABEL</type>
<position>-40,-13.5</position>
<gparam>LABEL_TEXT Set p/r</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1161</ID>
<type>DE_TO</type>
<position>-31.5,-20</position>
<input>
<ID>IN_0</ID>1284 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>1164</ID>
<type>DA_FROM</type>
<position>-58.5,-21</position>
<input>
<ID>IN_0</ID>1283 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>1166</ID>
<type>DA_FROM</type>
<position>-58.5,-23</position>
<input>
<ID>IN_0</ID>1282 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T3</lparam></gate>
<gate>
<ID>1174</ID>
<type>AA_AND2</type>
<position>-53.5,-22</position>
<input>
<ID>IN_0</ID>1283 </input>
<input>
<ID>IN_1</ID>1282 </input>
<output>
<ID>OUT</ID>1287 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1179</ID>
<type>DE_TO</type>
<position>-31.5,-24</position>
<input>
<ID>IN_0</ID>1289 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>15</ID>
<type>FF_GND</type>
<position>161.5,-108.5</position>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1182</ID>
<type>AA_LABEL</type>
<position>-40,-30.5</position>
<gparam>LABEL_TEXT Set DR_zero/AC_zero</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1189</ID>
<type>DE_TO</type>
<position>-31.5,-41.5</position>
<input>
<ID>IN_0</ID>1296 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR_zero</lparam></gate>
<gate>
<ID>1190</ID>
<type>AA_AND2</type>
<position>-36.5,-59</position>
<input>
<ID>IN_0</ID>1017 </input>
<input>
<ID>IN_1</ID>1018 </input>
<output>
<ID>OUT</ID>1299 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>AE_OR2</type>
<position>129,-215</position>
<input>
<ID>IN_0</ID>333 </input>
<input>
<ID>IN_1</ID>344 </input>
<output>
<ID>OUT</ID>153 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1193</ID>
<type>DE_TO</type>
<position>-31.5,-59</position>
<input>
<ID>IN_0</ID>1299 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC_zero</lparam></gate>
<gate>
<ID>1195</ID>
<type>DA_FROM</type>
<position>-56,-35</position>
<input>
<ID>IN_0</ID>360 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr1</lparam></gate>
<gate>
<ID>1196</ID>
<type>DA_FROM</type>
<position>-48.5,-36</position>
<input>
<ID>IN_0</ID>358 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr2</lparam></gate>
<gate>
<ID>1200</ID>
<type>DA_FROM</type>
<position>-48.5,-40</position>
<input>
<ID>IN_0</ID>359 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr6</lparam></gate>
<gate>
<ID>1201</ID>
<type>DA_FROM</type>
<position>-56,-41</position>
<input>
<ID>IN_0</ID>363 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr7</lparam></gate>
<gate>
<ID>1206</ID>
<type>DA_FROM</type>
<position>-48.5,-46</position>
<input>
<ID>IN_0</ID>384 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr12</lparam></gate>
<gate>
<ID>1207</ID>
<type>DA_FROM</type>
<position>-56,-47</position>
<input>
<ID>IN_0</ID>387 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr13</lparam></gate>
<gate>
<ID>1209</ID>
<type>DA_FROM</type>
<position>-56,-49</position>
<input>
<ID>IN_0</ID>388 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID dr15</lparam></gate>
<gate>
<ID>1224</ID>
<type>DA_FROM</type>
<position>-56,-52.5</position>
<input>
<ID>IN_0</ID>394 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac1</lparam></gate>
<gate>
<ID>1225</ID>
<type>DA_FROM</type>
<position>-48.5,-53.5</position>
<input>
<ID>IN_0</ID>392 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac2</lparam></gate>
<gate>
<ID>1227</ID>
<type>DA_FROM</type>
<position>-48.5,-55.5</position>
<input>
<ID>IN_0</ID>393 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac4</lparam></gate>
<gate>
<ID>1230</ID>
<type>DA_FROM</type>
<position>-56,-58.5</position>
<input>
<ID>IN_0</ID>431 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac7</lparam></gate>
<gate>
<ID>1232</ID>
<type>DA_FROM</type>
<position>-56,-60.5</position>
<input>
<ID>IN_0</ID>567 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac9</lparam></gate>
<gate>
<ID>1233</ID>
<type>DA_FROM</type>
<position>-48.5,-61.5</position>
<input>
<ID>IN_0</ID>539 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac10</lparam></gate>
<gate>
<ID>1235</ID>
<type>DA_FROM</type>
<position>-48.5,-63.5</position>
<input>
<ID>IN_0</ID>552 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac12</lparam></gate>
<gate>
<ID>1236</ID>
<type>DA_FROM</type>
<position>-56,-64.5</position>
<input>
<ID>IN_0</ID>598 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac13</lparam></gate>
<gate>
<ID>1238</ID>
<type>DA_FROM</type>
<position>-56,-66.5</position>
<input>
<ID>IN_0</ID>752 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ac15</lparam></gate>
<gate>
<ID>1239</ID>
<type>AA_LABEL</type>
<position>-42,-1.5</position>
<gparam>LABEL_TEXT Set</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>1240</ID>
<type>AA_LABEL</type>
<position>-40,-74</position>
<gparam>LABEL_TEXT Set AND/ADD/DR/INPR/COM/SHR/SHL</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1243</ID>
<type>DE_TO</type>
<position>-38,-90.5</position>
<input>
<ID>IN_0</ID>1346 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR</lparam></gate>
<gate>
<ID>1246</ID>
<type>DE_TO</type>
<position>-38,-108</position>
<input>
<ID>IN_0</ID>1355 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SHR</lparam></gate>
<gate>
<ID>1250</ID>
<type>DA_FROM</type>
<position>-48,-79.5</position>
<input>
<ID>IN_0</ID>1341 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>1284</ID>
<type>DA_FROM</type>
<position>-44.5,-144</position>
<input>
<ID>IN_0</ID>1369 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir8</lparam></gate>
<gate>
<ID>1251</ID>
<type>DA_FROM</type>
<position>-48,-81.5</position>
<input>
<ID>IN_0</ID>1342 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>1254</ID>
<type>DA_FROM</type>
<position>-48,-85</position>
<input>
<ID>IN_0</ID>1343 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>1256</ID>
<type>DA_FROM</type>
<position>-48,-90.5</position>
<input>
<ID>IN_0</ID>1346 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>1282</ID>
<type>DA_FROM</type>
<position>-44.5,-140</position>
<input>
<ID>IN_0</ID>1367 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir6</lparam></gate>
<gate>
<ID>1257</ID>
<type>DA_FROM</type>
<position>-48,-96</position>
<input>
<ID>IN_0</ID>1348 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B11</lparam></gate>
<gate>
<ID>1292</ID>
<type>DE_TO</type>
<position>-40.5,-134</position>
<input>
<ID>IN_0</ID>1364 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B3</lparam></gate>
<gate>
<ID>1259</ID>
<type>DA_FROM</type>
<position>-48,-94</position>
<input>
<ID>IN_0</ID>1347 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>1286</ID>
<type>DA_FROM</type>
<position>-44.5,-148</position>
<input>
<ID>IN_0</ID>1371 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir10</lparam></gate>
<gate>
<ID>1261</ID>
<type>AE_OR2</type>
<position>-49,-100.5</position>
<input>
<ID>IN_0</ID>1350 </input>
<input>
<ID>IN_1</ID>1351 </input>
<output>
<ID>OUT</ID>1353 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1262</ID>
<type>DA_FROM</type>
<position>-54,-99.5</position>
<input>
<ID>IN_0</ID>1350 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B8</lparam></gate>
<gate>
<ID>1280</ID>
<type>DA_FROM</type>
<position>-44.5,-136</position>
<input>
<ID>IN_0</ID>1365 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir4</lparam></gate>
<gate>
<ID>1263</ID>
<type>DA_FROM</type>
<position>-54,-101.5</position>
<input>
<ID>IN_0</ID>1351 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B9</lparam></gate>
<gate>
<ID>422</ID>
<type>DA_FROM</type>
<position>107.5,-88</position>
<input>
<ID>IN_0</ID>596 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID START</lparam></gate>
<gate>
<ID>1290</ID>
<type>DE_TO</type>
<position>-40.5,-130</position>
<input>
<ID>IN_0</ID>1362 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B1</lparam></gate>
<gate>
<ID>1265</ID>
<type>AA_AND2</type>
<position>-43,-101.5</position>
<input>
<ID>IN_0</ID>1353 </input>
<input>
<ID>IN_1</ID>1354 </input>
<output>
<ID>OUT</ID>1352 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1270</ID>
<type>DA_FROM</type>
<position>-48,-109</position>
<input>
<ID>IN_0</ID>1357 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B7</lparam></gate>
<gate>
<ID>1298</ID>
<type>DE_TO</type>
<position>-40.5,-146</position>
<input>
<ID>IN_0</ID>1370 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B9</lparam></gate>
<gate>
<ID>1273</ID>
<type>DA_FROM</type>
<position>-48,-115</position>
<input>
<ID>IN_0</ID>1359 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B6</lparam></gate>
<gate>
<ID>1274</ID>
<type>AA_LABEL</type>
<position>-42.5,-123</position>
<gparam>LABEL_TEXT Set B[i]</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1277</ID>
<type>DA_FROM</type>
<position>-44.5,-130</position>
<input>
<ID>IN_0</ID>1362 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir1</lparam></gate>
<gate>
<ID>1278</ID>
<type>DA_FROM</type>
<position>-44.5,-132</position>
<input>
<ID>IN_0</ID>1363 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir2</lparam></gate>
<gate>
<ID>1296</ID>
<type>DE_TO</type>
<position>-40.5,-142</position>
<input>
<ID>IN_0</ID>1368 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B7</lparam></gate>
<gate>
<ID>1279</ID>
<type>DA_FROM</type>
<position>-44.5,-134</position>
<input>
<ID>IN_0</ID>1364 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir3</lparam></gate>
<gate>
<ID>1287</ID>
<type>DA_FROM</type>
<position>-44.5,-150</position>
<input>
<ID>IN_0</ID>1372 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ir11</lparam></gate>
<gate>
<ID>1289</ID>
<type>DE_TO</type>
<position>-40.5,-128</position>
<input>
<ID>IN_0</ID>1361 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B0</lparam></gate>
<gate>
<ID>241</ID>
<type>DA_FROM</type>
<position>262.5,-23.5</position>
<input>
<ID>IN_0</ID>343 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>284</ID>
<type>CC_PULSE</type>
<position>250.5,-28.5</position>
<output>
<ID>OUT_0</ID>576 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 40</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>293</ID>
<type>DE_TO</type>
<position>264,-17</position>
<input>
<ID>IN_0</ID>560 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID START</lparam></gate>
<gate>
<ID>322</ID>
<type>DA_FROM</type>
<position>261,-39</position>
<input>
<ID>IN_0</ID>569 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID S</lparam></gate>
<gate>
<ID>339</ID>
<type>DA_FROM</type>
<position>261,-41</position>
<input>
<ID>IN_0</ID>572 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID START</lparam></gate>
<gate>
<ID>346</ID>
<type>AE_OR2</type>
<position>255.5,-25.5</position>
<input>
<ID>IN_0</ID>584 </input>
<input>
<ID>IN_1</ID>576 </input>
<output>
<ID>OUT</ID>586 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>363</ID>
<type>AA_LABEL</type>
<position>253,-19</position>
<gparam>LABEL_TEXT MANUAL START</gparam>
<gparam>TEXT_HEIGHT 0.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>431</ID>
<type>AA_LABEL</type>
<position>266.5,-30.5</position>
<gparam>LABEL_TEXT Clock</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>439</ID>
<type>AA_LABEL</type>
<position>265,-14.5</position>
<gparam>LABEL_TEXT Switch pulses are 2x the clock half-period</gparam>
<gparam>TEXT_HEIGHT 0.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>153</ID>
<type>DA_FROM</type>
<position>16,-67</position>
<input>
<ID>IN_0</ID>349 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>313</ID>
<type>DM_NOR8</type>
<position>-43.5,-55</position>
<input>
<ID>IN_0</ID>391 </input>
<input>
<ID>IN_1</ID>394 </input>
<input>
<ID>IN_2</ID>392 </input>
<input>
<ID>IN_3</ID>395 </input>
<input>
<ID>IN_4</ID>431 </input>
<input>
<ID>IN_5</ID>390 </input>
<input>
<ID>IN_6</ID>428 </input>
<input>
<ID>IN_7</ID>393 </input>
<output>
<ID>OUT</ID>1017 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>325</ID>
<type>DM_NOR8</type>
<position>-43.5,-63</position>
<input>
<ID>IN_0</ID>538 </input>
<input>
<ID>IN_1</ID>567 </input>
<input>
<ID>IN_2</ID>539 </input>
<input>
<ID>IN_3</ID>589 </input>
<input>
<ID>IN_4</ID>752 </input>
<input>
<ID>IN_5</ID>562 </input>
<input>
<ID>IN_6</ID>598 </input>
<input>
<ID>IN_7</ID>552 </input>
<output>
<ID>OUT</ID>1018 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<wire>
<ID>1122 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>217.5,-29.5,217.5,-29.5</points>
<connection>
<GID>957</GID>
<name>IN_0</name></connection>
<connection>
<GID>968</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>357 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46.5,-34,-46.5,-34</points>
<connection>
<GID>275</GID>
<name>IN_0</name></connection>
<connection>
<GID>1194</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>692 </ID>
<shape>
<vsegment>
<ID>4</ID>
<points>-112,-20.5,-112,-19.5</points>
<connection>
<GID>389</GID>
<name>ENABLE</name></connection>
<connection>
<GID>426</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1146 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>237.5,-57,237.5,-57</points>
<connection>
<GID>1005</GID>
<name>IN_0</name></connection>
<connection>
<GID>1003</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>150 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246.5,-25.5,246.5,-25.5</points>
<connection>
<GID>140</GID>
<name>IN_1</name></connection>
<connection>
<GID>1017</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1043 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>192,-85,192,-85</points>
<connection>
<GID>845</GID>
<name>OUT</name></connection>
<connection>
<GID>827</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>713 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150.5,-18,150.5,-18</points>
<connection>
<GID>451</GID>
<name>IN_0</name></connection>
<connection>
<GID>490</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>665 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-112,-25.5,-112,-25.5</points>
<connection>
<GID>389</GID>
<name>IN_2</name></connection>
<connection>
<GID>396</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1348 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46,-96,-46,-96</points>
<connection>
<GID>1258</GID>
<name>IN_1</name></connection>
<connection>
<GID>1257</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>151 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246.5,-23.5,246.5,-23.5</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<connection>
<GID>1016</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>345 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>180,-84,186,-84</points>
<connection>
<GID>845</GID>
<name>IN_0</name></connection>
<connection>
<GID>832</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>680 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-106,-27.5,-106,-27.5</points>
<connection>
<GID>389</GID>
<name>OUT_0</name></connection>
<connection>
<GID>400</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1134 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>228.5,-19.5,233.5,-19.5</points>
<connection>
<GID>967</GID>
<name>IN_0</name></connection>
<connection>
<GID>969</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>648 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-19,108.5,-14</points>
<connection>
<GID>374</GID>
<name>OUT</name></connection>
<connection>
<GID>387</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1070 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-172,111.5,-172</points>
<connection>
<GID>878</GID>
<name>IN_0</name></connection>
<connection>
<GID>879</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>584 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>252.5,-24.5,252.5,-24.5</points>
<connection>
<GID>140</GID>
<name>OUT</name></connection>
<connection>
<GID>346</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1237 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-114.5,29.5,-114.5</points>
<connection>
<GID>1113</GID>
<name>IN_0</name></connection>
<connection>
<GID>1114</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1109 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155.5,-215,155.5,-215</points>
<connection>
<GID>935</GID>
<name>OUT</name></connection>
<connection>
<GID>932</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>776 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,-56,125.5,-56</points>
<connection>
<GID>555</GID>
<name>IN_0</name></connection>
<connection>
<GID>572</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>759 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97,-55,97,-51.5</points>
<connection>
<GID>544</GID>
<name>OUT</name></connection>
<connection>
<GID>553</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1045 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186,-88.5,186,-86</points>
<connection>
<GID>843</GID>
<name>OUT</name></connection>
<connection>
<GID>845</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>615 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98.5,-19,98.5,-19</points>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<connection>
<GID>319</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1352 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40,-101.5,-40,-101.5</points>
<connection>
<GID>1245</GID>
<name>IN_0</name></connection>
<connection>
<GID>1265</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>814 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81.5,-86.5,81.5,-85.5</points>
<connection>
<GID>697</GID>
<name>OUT</name></connection>
<intersection>-85.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>81.5,-85.5,82,-85.5</points>
<connection>
<GID>757</GID>
<name>IN_1</name></connection>
<intersection>81.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>661 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-112,-27.5,-112,-27.5</points>
<connection>
<GID>389</GID>
<name>IN_0</name></connection>
<connection>
<GID>391</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1269 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-132,45,-132</points>
<connection>
<GID>1154</GID>
<name>IN_0</name></connection>
<connection>
<GID>1150</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1141 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>237.5,-48.5,237.5,-48.5</points>
<connection>
<GID>997</GID>
<name>OUT</name></connection>
<connection>
<GID>999</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>663 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-118.5,-26.5,-112,-26.5</points>
<connection>
<GID>389</GID>
<name>IN_1</name></connection>
<connection>
<GID>393</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>687 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-106,-26.5,-101,-26.5</points>
<connection>
<GID>389</GID>
<name>OUT_1</name></connection>
<connection>
<GID>410</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>670 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-106,-25.5,-106,-25.5</points>
<connection>
<GID>389</GID>
<name>OUT_2</name></connection>
<connection>
<GID>398</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1231 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-104.5,37,-104.5</points>
<connection>
<GID>1106</GID>
<name>IN_0</name></connection>
<connection>
<GID>1108</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>685 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-106,-24.5,-101,-24.5</points>
<connection>
<GID>389</GID>
<name>OUT_3</name></connection>
<connection>
<GID>411</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>827 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>103.5,-85,103.5,-85</points>
<connection>
<GID>761</GID>
<name>IN_0</name></connection>
<connection>
<GID>762</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1034 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>159.5,-102,161.5,-102</points>
<connection>
<GID>818</GID>
<name>IN_3</name></connection>
<intersection>159.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>159.5,-106,159.5,-102</points>
<intersection>-106 11</intersection>
<intersection>-102 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>145.5,-106,159.5,-106</points>
<connection>
<GID>805</GID>
<name>OUT</name></connection>
<intersection>159.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>333 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126,-214,126,-214</points>
<connection>
<GID>929</GID>
<name>OUT</name></connection>
<connection>
<GID>10</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>668 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-106,-23.5,-106,-23.5</points>
<connection>
<GID>389</GID>
<name>OUT_4</name></connection>
<connection>
<GID>413</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>683 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-106,-22.5,-101,-22.5</points>
<connection>
<GID>389</GID>
<name>OUT_5</name></connection>
<connection>
<GID>415</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1030 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133.5,-126.5,133.5,-124.5</points>
<connection>
<GID>826</GID>
<name>IN_1</name></connection>
<connection>
<GID>812</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>672 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-106,-21.5,-106,-21.5</points>
<connection>
<GID>389</GID>
<name>OUT_6</name></connection>
<connection>
<GID>417</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1371 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,-148,-42.5,-148</points>
<connection>
<GID>1299</GID>
<name>IN_0</name></connection>
<connection>
<GID>1286</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>682 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-106,-20.5,-101,-20.5</points>
<connection>
<GID>389</GID>
<name>OUT_7</name></connection>
<connection>
<GID>419</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>644 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-19,102.5,-19</points>
<connection>
<GID>319</GID>
<name>OUT_0</name></connection>
<connection>
<GID>377</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1266 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-130,51,-130</points>
<connection>
<GID>1151</GID>
<name>IN_0</name></connection>
<connection>
<GID>1149</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>1074 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-172,141.5,-172</points>
<connection>
<GID>883</GID>
<name>IN_0</name></connection>
<connection>
<GID>882</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1140 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230.5,-51.5,230.5,-51.5</points>
<connection>
<GID>991</GID>
<name>IN_0</name></connection>
<connection>
<GID>997</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>1076 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145.5,-172,145.5,-172</points>
<connection>
<GID>883</GID>
<name>OUT_0</name></connection>
<connection>
<GID>885</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>428 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-54,-56.5,-46.5,-56.5</points>
<connection>
<GID>313</GID>
<name>IN_6</name></connection>
<connection>
<GID>1228</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1296 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33.5,-41.5,-33.5,-41.5</points>
<connection>
<GID>1188</GID>
<name>OUT</name></connection>
<connection>
<GID>1189</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1360 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40,-114,-40,-114</points>
<connection>
<GID>1247</GID>
<name>IN_0</name></connection>
<connection>
<GID>1271</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>761 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97,-61,97,-57</points>
<connection>
<GID>553</GID>
<name>IN_1</name></connection>
<intersection>-61 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>96.5,-61,97,-61</points>
<connection>
<GID>548</GID>
<name>OUT</name></connection>
<intersection>97 0</intersection></hsegment></shape></wire>
<wire>
<ID>757 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,-56,103,-56</points>
<connection>
<GID>553</GID>
<name>OUT</name></connection>
<connection>
<GID>505</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>792 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>172,-55,172,-54</points>
<connection>
<GID>597</GID>
<name>OUT</name></connection>
<intersection>-55 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>172,-55,172.5,-55</points>
<connection>
<GID>615</GID>
<name>IN_0</name></connection>
<intersection>172 0</intersection></hsegment></shape></wire>
<wire>
<ID>1125 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222.5,-26.5,222.5,-26.5</points>
<connection>
<GID>968</GID>
<name>OUT_0</name></connection>
<connection>
<GID>969</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1342 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46,-81.5,-46,-81.5</points>
<connection>
<GID>1249</GID>
<name>IN_1</name></connection>
<connection>
<GID>1251</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>711 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150.5,-16,150.5,-16</points>
<connection>
<GID>448</GID>
<name>IN_0</name></connection>
<connection>
<GID>490</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>709 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150.5,-25,150.5,-24</points>
<connection>
<GID>480</GID>
<name>IN_1</name></connection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>144.5,-25,150.5,-25</points>
<connection>
<GID>468</GID>
<name>IN_0</name></connection>
<intersection>150.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1131 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228.5,-22.5,228.5,-22.5</points>
<connection>
<GID>964</GID>
<name>IN_0</name></connection>
<connection>
<GID>969</GID>
<name>OUT_4</name></connection></vsegment></shape></wire>
<wire>
<ID>641 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-23,102.5,-23</points>
<connection>
<GID>334</GID>
<name>IN_0</name></connection>
<connection>
<GID>377</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>1340 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40,-80.5,-40,-80.5</points>
<connection>
<GID>1241</GID>
<name>IN_0</name></connection>
<connection>
<GID>1249</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>1136 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219.5,-29.5,219.5,-29.5</points>
<connection>
<GID>968</GID>
<name>clear</name></connection>
<connection>
<GID>958</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1086 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-192,115.5,-192</points>
<connection>
<GID>890</GID>
<name>IN_0</name></connection>
<connection>
<GID>893</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>600 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>218.5,-20.5,219.5,-20.5</points>
<connection>
<GID>955</GID>
<name>OUT_0</name></connection>
<connection>
<GID>968</GID>
<name>count_enable</name></connection>
<connection>
<GID>968</GID>
<name>count_up</name></connection></hsegment></shape></wire>
<wire>
<ID>1126 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222.5,-25.5,222.5,-25.5</points>
<connection>
<GID>968</GID>
<name>OUT_1</name></connection>
<connection>
<GID>969</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1347 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46,-94,-46,-94</points>
<connection>
<GID>1258</GID>
<name>IN_0</name></connection>
<connection>
<GID>1259</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>658 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-21,108.5,-21</points>
<connection>
<GID>387</GID>
<name>IN_1</name></connection>
<connection>
<GID>377</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>1124 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222.5,-24.5,222.5,-24.5</points>
<connection>
<GID>968</GID>
<name>OUT_2</name></connection>
<connection>
<GID>969</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>831 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-81.5,135.5,-81.5</points>
<connection>
<GID>766</GID>
<name>IN_0</name></connection>
<connection>
<GID>764</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>613 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98.5,-13,98.5,-13</points>
<connection>
<GID>296</GID>
<name>IN_0</name></connection>
<connection>
<GID>300</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1022 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139.5,-81.5,139.5,-81.5</points>
<connection>
<GID>766</GID>
<name>OUT_0</name></connection>
<connection>
<GID>820</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>646 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-21,114.5,-21</points>
<connection>
<GID>289</GID>
<name>IN_0</name></connection>
<connection>
<GID>387</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>1005 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139.5,-105,139.5,-105</points>
<connection>
<GID>805</GID>
<name>IN_0</name></connection>
<connection>
<GID>808</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>1025 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139.5,-89,139.5,-89</points>
<connection>
<GID>769</GID>
<name>IN_0</name></connection>
<connection>
<GID>822</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1004 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139.5,-117,139.5,-107</points>
<connection>
<GID>805</GID>
<name>IN_1</name></connection>
<intersection>-117 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>125.5,-117,139.5,-117</points>
<connection>
<GID>781</GID>
<name>IN_0</name></connection>
<intersection>139.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>359 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46.5,-40,-46.5,-40</points>
<connection>
<GID>275</GID>
<name>IN_5</name></connection>
<connection>
<GID>1200</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>706 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144.5,-23,144.5,-23</points>
<connection>
<GID>467</GID>
<name>IN_0</name></connection>
<connection>
<GID>476</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>560 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>257,-21.5,264.5,-21.5</points>
<connection>
<GID>18</GID>
<name>J</name></connection>
<connection>
<GID>285</GID>
<name>OUT_0</name></connection>
<intersection>257 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>257,-21.5,257,-17</points>
<intersection>-21.5 1</intersection>
<intersection>-17 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>257,-17,262,-17</points>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<intersection>257 7</intersection></hsegment></shape></wire>
<wire>
<ID>1135 </ID>
<shape>
<vsegment>
<ID>11</ID>
<points>222.5,-19.5,222.5,-18.5</points>
<connection>
<GID>969</GID>
<name>ENABLE</name></connection>
<connection>
<GID>971</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1008 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,-110,132,-106</points>
<intersection>-110 2</intersection>
<intersection>-106 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132,-106,132.5,-106</points>
<connection>
<GID>808</GID>
<name>IN_2</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>131.5,-110,132,-110</points>
<connection>
<GID>799</GID>
<name>OUT</name></connection>
<intersection>132 0</intersection></hsegment></shape></wire>
<wire>
<ID>1366 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,-138,-42.5,-138</points>
<connection>
<GID>1281</GID>
<name>IN_0</name></connection>
<connection>
<GID>1294</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1234 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-112.5,29.5,-112.5</points>
<connection>
<GID>1110</GID>
<name>IN_0</name></connection>
<connection>
<GID>1112</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>637 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-13,102.5,-13</points>
<connection>
<GID>300</GID>
<name>OUT_0</name></connection>
<connection>
<GID>374</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1354 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46,-103.5,-46,-102.5</points>
<connection>
<GID>1265</GID>
<name>IN_1</name></connection>
<intersection>-103.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-52,-103.5,-46,-103.5</points>
<connection>
<GID>1266</GID>
<name>IN_0</name></connection>
<intersection>-46 0</intersection></hsegment></shape></wire>
<wire>
<ID>635 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-15,102.5,-15</points>
<connection>
<GID>311</GID>
<name>IN_0</name></connection>
<connection>
<GID>374</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>639 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-21,102.5,-21</points>
<connection>
<GID>323</GID>
<name>IN_0</name></connection>
<connection>
<GID>377</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1012 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127.5,-123.5,127.5,-123.5</points>
<connection>
<GID>789</GID>
<name>IN_0</name></connection>
<connection>
<GID>810</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>659 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-29.5,108.5,-23</points>
<connection>
<GID>369</GID>
<name>OUT</name></connection>
<connection>
<GID>387</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>1169 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-44,18,-44</points>
<connection>
<GID>1030</GID>
<name>IN_0</name></connection>
<connection>
<GID>1040</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>617 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>89.5,-25.5,95.5,-25.5</points>
<connection>
<GID>337</GID>
<name>IN_0</name></connection>
<connection>
<GID>365</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1166 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-38,18,-38</points>
<connection>
<GID>1028</GID>
<name>IN_0</name></connection>
<connection>
<GID>1039</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>620 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>89.5,-27.5,95.5,-27.5</points>
<connection>
<GID>343</GID>
<name>IN_0</name></connection>
<connection>
<GID>365</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>622 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>89.5,-29.5,95.5,-29.5</points>
<connection>
<GID>348</GID>
<name>IN_0</name></connection>
<connection>
<GID>365</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1010 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,-113,125.5,-113</points>
<connection>
<GID>806</GID>
<name>IN_0</name></connection>
<connection>
<GID>784</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1011 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,-115,125.5,-115</points>
<connection>
<GID>806</GID>
<name>IN_1</name></connection>
<connection>
<GID>785</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1009 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,-114,132.5,-108</points>
<connection>
<GID>808</GID>
<name>IN_3</name></connection>
<intersection>-114 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>131.5,-114,132.5,-114</points>
<connection>
<GID>806</GID>
<name>OUT</name></connection>
<intersection>132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>704 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144.5,-21,144.5,-21</points>
<connection>
<GID>476</GID>
<name>IN_0</name></connection>
<connection>
<GID>455</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>707 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150.5,-22,150.5,-22</points>
<connection>
<GID>476</GID>
<name>OUT</name></connection>
<connection>
<GID>480</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>624 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>89.5,-31.5,95.5,-31.5</points>
<connection>
<GID>351</GID>
<name>IN_0</name></connection>
<connection>
<GID>365</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1225 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-91,40.5,-91</points>
<connection>
<GID>1100</GID>
<name>IN_0</name></connection>
<connection>
<GID>1098</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1224 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-93,40.5,-93</points>
<connection>
<GID>1100</GID>
<name>IN_1</name></connection>
<connection>
<GID>1097</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1227 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-92,46.5,-89</points>
<connection>
<GID>1058</GID>
<name>K</name></connection>
<connection>
<GID>1100</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>634 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-33.5,102.5,-30.5</points>
<connection>
<GID>369</GID>
<name>IN_1</name></connection>
<intersection>-33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89.5,-33.5,102.5,-33.5</points>
<connection>
<GID>362</GID>
<name>IN_0</name></connection>
<intersection>102.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1144 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>231.5,-56,231.5,-56</points>
<connection>
<GID>1003</GID>
<name>IN_0</name></connection>
<connection>
<GID>986</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>148 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,-59,86.5,-59</points>
<connection>
<GID>527</GID>
<name>IN_0</name></connection>
<connection>
<GID>1</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>383 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46.5,-42,-46.5,-42</points>
<connection>
<GID>1202</GID>
<name>IN_0</name></connection>
<connection>
<GID>287</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1068 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163,-152,163,-150</points>
<connection>
<GID>875</GID>
<name>OUT</name></connection>
<connection>
<GID>872</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>730 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-21,156.5,-17</points>
<connection>
<GID>498</GID>
<name>IN_0</name></connection>
<connection>
<GID>490</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>1349 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40,-95,-40,-95</points>
<connection>
<GID>1258</GID>
<name>OUT</name></connection>
<connection>
<GID>1244</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>632 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-28.5,102.5,-28.5</points>
<connection>
<GID>365</GID>
<name>OUT</name></connection>
<connection>
<GID>369</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1197 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-87,46.5,-87</points>
<connection>
<GID>1062</GID>
<name>IN_0</name></connection>
<connection>
<GID>1058</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>1083 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145.5,-194,145.5,-194</points>
<connection>
<GID>895</GID>
<name>IN_0</name></connection>
<connection>
<GID>896</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>778 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>143,-55,143,-55</points>
<connection>
<GID>576</GID>
<name>IN_0</name></connection>
<connection>
<GID>581</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>586 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>258.5,-25.5,264.5,-25.5</points>
<connection>
<GID>18</GID>
<name>K</name></connection>
<connection>
<GID>346</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1028 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133.5,-122.5,133.5,-122.5</points>
<connection>
<GID>810</GID>
<name>OUT</name></connection>
<connection>
<GID>826</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>343 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>264.5,-23.5,264.5,-23.5</points>
<connection>
<GID>18</GID>
<name>clock</name></connection>
<connection>
<GID>241</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>785 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,-55,166,-55</points>
<connection>
<GID>594</GID>
<name>IN_0</name></connection>
<connection>
<GID>597</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>96 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>270.5,-21.5,270.5,-21.5</points>
<connection>
<GID>18</GID>
<name>Q</name></connection>
<connection>
<GID>1013</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1200 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-85.5,22.5,-85.5</points>
<connection>
<GID>1070</GID>
<name>IN_0</name></connection>
<connection>
<GID>1066</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1221 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-85.5,27,-83.5</points>
<intersection>-85.5 2</intersection>
<intersection>-83.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-85.5,27,-85.5</points>
<connection>
<GID>1070</GID>
<name>OUT_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>27,-83.5,29,-83.5</points>
<connection>
<GID>1096</GID>
<name>IN_2</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>1153 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>243.5,-48.5,258.5,-48.5</points>
<connection>
<GID>1011</GID>
<name>IN_0</name></connection>
<intersection>243.5 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>243.5,-48.5,243.5,-42</points>
<connection>
<GID>1007</GID>
<name>OUT</name></connection>
<intersection>-48.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>1367 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,-140,-42.5,-140</points>
<connection>
<GID>1295</GID>
<name>IN_0</name></connection>
<connection>
<GID>1282</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>385 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-54,-43,-46.5,-43</points>
<connection>
<GID>1203</GID>
<name>IN_0</name></connection>
<connection>
<GID>287</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>720 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162.5,-23,162.5,-23</points>
<connection>
<GID>444</GID>
<name>IN_0</name></connection>
<connection>
<GID>498</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>716 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150.5,-29,150.5,-29</points>
<connection>
<GID>470</GID>
<name>IN_0</name></connection>
<connection>
<GID>494</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1149 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>237.5,-41,237.5,-41</points>
<connection>
<GID>975</GID>
<name>IN_0</name></connection>
<connection>
<GID>1007</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>816 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-84.5,88,-84.5</points>
<connection>
<GID>619</GID>
<name>IN_0</name></connection>
<connection>
<GID>757</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>355 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-68,27.5,-65</points>
<intersection>-68 2</intersection>
<intersection>-65 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-65,31.5,-65</points>
<connection>
<GID>249</GID>
<name>IN_3</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-68,27.5,-68</points>
<connection>
<GID>39</GID>
<name>OUT</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>718 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150.5,-27,150.5,-27</points>
<connection>
<GID>472</GID>
<name>IN_0</name></connection>
<connection>
<GID>494</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>393 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46.5,-55.5,-46.5,-55.5</points>
<connection>
<GID>1227</GID>
<name>IN_0</name></connection>
<connection>
<GID>313</GID>
<name>IN_7</name></connection></vsegment></shape></wire>
<wire>
<ID>728 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-23,156.5,-23</points>
<connection>
<GID>480</GID>
<name>OUT</name></connection>
<connection>
<GID>498</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1013 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127.5,-121.5,127.5,-121.5</points>
<connection>
<GID>810</GID>
<name>IN_0</name></connection>
<connection>
<GID>788</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>731 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-28,156.5,-25</points>
<connection>
<GID>498</GID>
<name>IN_2</name></connection>
<connection>
<GID>494</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>733 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-49.5,81,-49.5</points>
<connection>
<GID>515</GID>
<name>IN_0</name></connection>
<connection>
<GID>516</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1102 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96,-222.5,96,-216.5</points>
<connection>
<GID>926</GID>
<name>IN_2</name></connection>
<connection>
<GID>924</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>744 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-50.5,91,-49.5</points>
<connection>
<GID>544</GID>
<name>IN_0</name></connection>
<intersection>-49.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>85,-49.5,91,-49.5</points>
<connection>
<GID>516</GID>
<name>OUT_0</name></connection>
<intersection>91 0</intersection></hsegment></shape></wire>
<wire>
<ID>1158 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245,-69,245,-53.5</points>
<intersection>-69 2</intersection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>245,-53.5,258.5,-53.5</points>
<connection>
<GID>1011</GID>
<name>IN_6</name></connection>
<intersection>245 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>243.5,-69,245,-69</points>
<connection>
<GID>995</GID>
<name>IN_0</name></connection>
<intersection>245 0</intersection></hsegment></shape></wire>
<wire>
<ID>740 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-51.5,85,-51.5</points>
<connection>
<GID>518</GID>
<name>IN_0</name></connection>
<connection>
<GID>540</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1147 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>237.5,-60,237.5,-59</points>
<connection>
<GID>1005</GID>
<name>IN_1</name></connection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>231.5,-60,237.5,-60</points>
<connection>
<GID>989</GID>
<name>IN_0</name></connection>
<intersection>237.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1155 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>243.5,-50.5,258.5,-50.5</points>
<connection>
<GID>1011</GID>
<name>IN_2</name></connection>
<intersection>243.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>243.5,-58,243.5,-50.5</points>
<connection>
<GID>1005</GID>
<name>OUT</name></connection>
<intersection>-50.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1267 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-128,51,-128</points>
<connection>
<GID>1149</GID>
<name>J</name></connection>
<connection>
<GID>1153</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>737 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-53.5,85,-53.5</points>
<connection>
<GID>524</GID>
<name>IN_0</name></connection>
<connection>
<GID>540</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1145 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>231.5,-58,231.5,-58</points>
<connection>
<GID>1003</GID>
<name>IN_1</name></connection>
<connection>
<GID>988</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1111 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>175.5,-218,175.5,-218</points>
<connection>
<GID>942</GID>
<name>IN_0</name></connection>
<connection>
<GID>943</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>565 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>264.5,-35.5,269,-35.5</points>
<connection>
<GID>317</GID>
<name>IN_0</name></connection>
<connection>
<GID>298</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>1112 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>175.5,-216,175.5,-216</points>
<connection>
<GID>941</GID>
<name>IN_0</name></connection>
<connection>
<GID>943</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>574 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269,-40,269,-37.5</points>
<connection>
<GID>335</GID>
<name>OUT</name></connection>
<connection>
<GID>317</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1282 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-56.5,-23,-56.5,-23</points>
<connection>
<GID>1166</GID>
<name>IN_0</name></connection>
<connection>
<GID>1174</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>563 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>275,-36.5,275,-36.5</points>
<connection>
<GID>317</GID>
<name>OUT</name></connection>
<connection>
<GID>310</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>788 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,-57,166,-57</points>
<connection>
<GID>599</GID>
<name>IN_0</name></connection>
<connection>
<GID>611</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>755 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-63,90.5,-63</points>
<connection>
<GID>528</GID>
<name>IN_0</name></connection>
<connection>
<GID>548</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>754 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-61,90.5,-61</points>
<connection>
<GID>530</GID>
<name>IN_0</name></connection>
<connection>
<GID>548</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>742 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-52.5,91,-52.5</points>
<connection>
<GID>540</GID>
<name>OUT</name></connection>
<connection>
<GID>544</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1243 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,-18.5,59,-18.5</points>
<connection>
<GID>1019</GID>
<name>IN_0</name></connection>
<connection>
<GID>1118</GID>
<name>Q</name></connection></vsegment></shape></wire>
<wire>
<ID>1185 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39,-44,50,-44</points>
<connection>
<GID>1037</GID>
<name>J</name></connection>
<intersection>39 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>39,-48.5,39,-44</points>
<connection>
<GID>1052</GID>
<name>IN_0</name></connection>
<connection>
<GID>1043</GID>
<name>OUT</name></connection>
<intersection>-44 1</intersection></vsegment></shape></wire>
<wire>
<ID>13 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-59,90.5,-59</points>
<connection>
<GID>548</GID>
<name>IN_0</name></connection>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>380 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-39.5,-40.5,-39.5,-37.5</points>
<connection>
<GID>1188</GID>
<name>IN_0</name></connection>
<connection>
<GID>275</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>1103 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-214.5,102,-214.5</points>
<connection>
<GID>899</GID>
<name>IN_0</name></connection>
<connection>
<GID>926</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>848 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,-101,125.5,-101</points>
<connection>
<GID>773</GID>
<name>OUT_0</name></connection>
<connection>
<GID>795</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1341 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46,-79.5,-46,-79.5</points>
<connection>
<GID>1249</GID>
<name>IN_0</name></connection>
<connection>
<GID>1250</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>766 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>119.5,-55,119.5,-55</points>
<connection>
<GID>567</GID>
<name>IN_0</name></connection>
<connection>
<GID>572</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>768 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>119.5,-57,119.5,-57</points>
<connection>
<GID>568</GID>
<name>IN_0</name></connection>
<connection>
<GID>572</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1107 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149.5,-214,149.5,-214</points>
<connection>
<GID>935</GID>
<name>IN_0</name></connection>
<connection>
<GID>936</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1108 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149.5,-216,149.5,-216</points>
<connection>
<GID>935</GID>
<name>IN_1</name></connection>
<connection>
<GID>937</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1370 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,-146,-42.5,-146</points>
<connection>
<GID>1285</GID>
<name>IN_0</name></connection>
<connection>
<GID>1298</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>781 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149,-56,149,-56</points>
<connection>
<GID>574</GID>
<name>IN_0</name></connection>
<connection>
<GID>581</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>539 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46.5,-61.5,-46.5,-61.5</points>
<connection>
<GID>325</GID>
<name>IN_2</name></connection>
<connection>
<GID>1233</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>390 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46.5,-57.5,-46.5,-57.5</points>
<connection>
<GID>1229</GID>
<name>IN_0</name></connection>
<connection>
<GID>313</GID>
<name>IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>1233 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-110.5,29.5,-110.5</points>
<connection>
<GID>1112</GID>
<name>IN_0</name></connection>
<connection>
<GID>1111</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>388 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-54,-49,-46.5,-49</points>
<connection>
<GID>287</GID>
<name>IN_4</name></connection>
<connection>
<GID>1209</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1239 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-113,36,-111.5</points>
<intersection>-113 1</intersection>
<intersection>-111.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-113,37,-113</points>
<connection>
<GID>1117</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-111.5,36,-111.5</points>
<connection>
<GID>1112</GID>
<name>OUT</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>1114 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>175.5,-214,175.5,-214</points>
<connection>
<GID>947</GID>
<name>IN_0</name></connection>
<connection>
<GID>948</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>779 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>143,-57,143,-57</points>
<connection>
<GID>579</GID>
<name>IN_0</name></connection>
<connection>
<GID>581</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1344 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46,-87,-46,-87</points>
<connection>
<GID>1255</GID>
<name>IN_0</name></connection>
<connection>
<GID>1253</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>802 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178.5,-56,178.5,-56</points>
<connection>
<GID>588</GID>
<name>IN_0</name></connection>
<connection>
<GID>615</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>783 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,-53,166,-53</points>
<connection>
<GID>591</GID>
<name>IN_0</name></connection>
<connection>
<GID>597</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1199 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-83.5,22.5,-83.5</points>
<connection>
<GID>1069</GID>
<name>IN_0</name></connection>
<connection>
<GID>1065</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>857 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,-111,125.5,-111</points>
<connection>
<GID>782</GID>
<name>IN_0</name></connection>
<connection>
<GID>799</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1220 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-83.5,26.5,-82.5</points>
<connection>
<GID>1069</GID>
<name>OUT_0</name></connection>
<intersection>-82.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-82.5,29,-82.5</points>
<connection>
<GID>1096</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1223 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-91,28,-85.5</points>
<intersection>-91 2</intersection>
<intersection>-85.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-85.5,29,-85.5</points>
<connection>
<GID>1096</GID>
<name>IN_4</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-91,28,-91</points>
<connection>
<GID>1076</GID>
<name>OUT</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>1368 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,-142,-42.5,-142</points>
<connection>
<GID>1283</GID>
<name>IN_0</name></connection>
<connection>
<GID>1296</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>153 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,-215,132,-215</points>
<connection>
<GID>927</GID>
<name>IN_0</name></connection>
<connection>
<GID>10</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>1358 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46,-113,-46,-113</points>
<connection>
<GID>1271</GID>
<name>IN_0</name></connection>
<connection>
<GID>1272</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1359 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46,-115,-46,-115</points>
<connection>
<GID>1271</GID>
<name>IN_1</name></connection>
<connection>
<GID>1273</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>790 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,-59,166,-59</points>
<connection>
<GID>601</GID>
<name>IN_0</name></connection>
<connection>
<GID>611</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1133 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228.5,-20.5,228.5,-20.5</points>
<connection>
<GID>966</GID>
<name>IN_0</name></connection>
<connection>
<GID>969</GID>
<name>OUT_6</name></connection></vsegment></shape></wire>
<wire>
<ID>800 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>172,-58,172,-57</points>
<connection>
<GID>611</GID>
<name>OUT</name></connection>
<intersection>-57 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>172,-57,172.5,-57</points>
<connection>
<GID>615</GID>
<name>IN_1</name></connection>
<intersection>172 0</intersection></hsegment></shape></wire>
<wire>
<ID>1138 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230.5,-45.5,230.5,-45.5</points>
<connection>
<GID>978</GID>
<name>IN_0</name></connection>
<connection>
<GID>997</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>803 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-81.5,75.5,-81.5</points>
<connection>
<GID>623</GID>
<name>IN_0</name></connection>
<connection>
<GID>626</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1351 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52,-101.5,-52,-101.5</points>
<connection>
<GID>1261</GID>
<name>IN_1</name></connection>
<connection>
<GID>1263</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>805 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-83.5,75.5,-83.5</points>
<connection>
<GID>625</GID>
<name>IN_0</name></connection>
<connection>
<GID>626</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>812 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81.5,-83.5,81.5,-82.5</points>
<connection>
<GID>626</GID>
<name>OUT</name></connection>
<intersection>-83.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>81.5,-83.5,82,-83.5</points>
<connection>
<GID>757</GID>
<name>IN_0</name></connection>
<intersection>81.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>807 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-85.5,75.5,-85.5</points>
<connection>
<GID>684</GID>
<name>IN_0</name></connection>
<connection>
<GID>697</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1172 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-52,18,-52</points>
<connection>
<GID>1034</GID>
<name>IN_0</name></connection>
<connection>
<GID>1041</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>809 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-87.5,75.5,-87.5</points>
<connection>
<GID>685</GID>
<name>IN_0</name></connection>
<connection>
<GID>697</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1069 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163,-148,163,-146</points>
<connection>
<GID>874</GID>
<name>OUT</name></connection>
<connection>
<GID>872</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>591 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-85,115.5,-85</points>
<connection>
<GID>758</GID>
<name>IN_0</name></connection>
<connection>
<GID>425</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>826 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>103.5,-83,103.5,-83</points>
<connection>
<GID>760</GID>
<name>IN_0</name></connection>
<connection>
<GID>762</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>572 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>263,-41,263,-41</points>
<connection>
<GID>335</GID>
<name>IN_1</name></connection>
<connection>
<GID>339</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1258 </ID>
<shape>
<vsegment>
<ID>5</ID>
<points>53,-18.5,53,-17.5</points>
<connection>
<GID>1118</GID>
<name>J</name></connection>
<intersection>-17.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>47,-17.5,53,-17.5</points>
<connection>
<GID>1125</GID>
<name>OUT</name></connection>
<intersection>53 5</intersection></hsegment></shape></wire>
<wire>
<ID>1273 </ID>
<shape>
<vsegment>
<ID>9</ID>
<points>53,-23.5,53,-22.5</points>
<connection>
<GID>1118</GID>
<name>K</name></connection>
<intersection>-23.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>47,-23.5,53,-23.5</points>
<connection>
<GID>1156</GID>
<name>OUT</name></connection>
<intersection>53 9</intersection></hsegment></shape></wire>
<wire>
<ID>1244 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-20.5,53,-20.5</points>
<connection>
<GID>1118</GID>
<name>clock</name></connection>
<connection>
<GID>1119</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>593 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-84,109.5,-84</points>
<connection>
<GID>425</GID>
<name>IN_0</name></connection>
<connection>
<GID>762</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>596 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-88,109.5,-86</points>
<connection>
<GID>422</GID>
<name>IN_0</name></connection>
<connection>
<GID>425</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1041 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>180,-89.5,180,-89.5</points>
<connection>
<GID>834</GID>
<name>IN_0</name></connection>
<connection>
<GID>843</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1020 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168.5,-102.5,168.5,-102.5</points>
<connection>
<GID>763</GID>
<name>IN_0</name></connection>
<connection>
<GID>818</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>1369 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,-144,-42.5,-144</points>
<connection>
<GID>1297</GID>
<name>IN_0</name></connection>
<connection>
<GID>1284</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1023 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139.5,-83.5,139.5,-83.5</points>
<connection>
<GID>767</GID>
<name>IN_0</name></connection>
<connection>
<GID>820</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>838 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-113,121.5,-113</points>
<connection>
<GID>784</GID>
<name>IN_0</name></connection>
<connection>
<GID>783</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1240 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-115.5,36,-115</points>
<intersection>-115.5 2</intersection>
<intersection>-115 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-115,37,-115</points>
<connection>
<GID>1117</GID>
<name>IN_1</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-115.5,36,-115.5</points>
<connection>
<GID>1114</GID>
<name>OUT</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>1242 </ID>
<shape>
<vsegment>
<ID>3</ID>
<points>43,-114,43,-112</points>
<connection>
<GID>1103</GID>
<name>K</name></connection>
<connection>
<GID>1117</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>1024 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139.5,-87,139.5,-87</points>
<connection>
<GID>768</GID>
<name>IN_0</name></connection>
<connection>
<GID>822</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1056 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>139.5,-96.5,139.5,-96.5</points>
<connection>
<GID>770</GID>
<name>IN_0</name></connection>
<connection>
<GID>864</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1057 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>139.5,-98.5,139.5,-98.5</points>
<connection>
<GID>771</GID>
<name>IN_0</name></connection>
<connection>
<GID>864</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1232 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-106.5,37,-106.5</points>
<connection>
<GID>1106</GID>
<name>IN_1</name></connection>
<connection>
<GID>1109</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1230 </ID>
<shape>
<vsegment>
<ID>4</ID>
<points>43,-108,43,-105.5</points>
<connection>
<GID>1103</GID>
<name>J</name></connection>
<connection>
<GID>1106</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>833 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-101,121.5,-101</points>
<connection>
<GID>772</GID>
<name>IN_0</name></connection>
<connection>
<GID>773</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1202 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-92,20.5,-92</points>
<connection>
<GID>1080</GID>
<name>IN_0</name></connection>
<connection>
<GID>1076</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>850 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,-103,125.5,-103</points>
<connection>
<GID>775</GID>
<name>IN_0</name></connection>
<connection>
<GID>795</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>851 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,-105,125.5,-105</points>
<connection>
<GID>776</GID>
<name>IN_0</name></connection>
<connection>
<GID>797</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>541 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>258.5,-56.5,258.5,-55.5</points>
<connection>
<GID>1011</GID>
<name>IN_4</name></connection>
<connection>
<GID>246</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1032 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,-100,160,-96</points>
<intersection>-100 1</intersection>
<intersection>-96 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>160,-100,161.5,-100</points>
<connection>
<GID>818</GID>
<name>IN_1</name></connection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>145.5,-96,160,-96</points>
<intersection>145.5 3</intersection>
<intersection>160 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>145.5,-96,145.5,-88</points>
<connection>
<GID>822</GID>
<name>OUT</name></connection>
<intersection>-96 2</intersection></vsegment></shape></wire>
<wire>
<ID>853 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,-107,125.5,-107</points>
<connection>
<GID>779</GID>
<name>IN_0</name></connection>
<connection>
<GID>797</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1238 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-116.5,29.5,-116.5</points>
<connection>
<GID>1114</GID>
<name>IN_1</name></connection>
<connection>
<GID>1115</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>855 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,-109,125.5,-109</points>
<connection>
<GID>780</GID>
<name>IN_0</name></connection>
<connection>
<GID>799</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1361 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,-128,-42.5,-128</points>
<connection>
<GID>1276</GID>
<name>IN_0</name></connection>
<connection>
<GID>1289</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1019 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>127.5,-125.5,139.5,-125.5</points>
<connection>
<GID>816</GID>
<name>IN_1</name></connection>
<intersection>127.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>127.5,-129.5,127.5,-125.5</points>
<connection>
<GID>790</GID>
<name>IN_0</name></connection>
<intersection>-125.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>1173 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-50,18,-50</points>
<connection>
<GID>1033</GID>
<name>IN_0</name></connection>
<connection>
<GID>1041</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>840 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123.5,-125.5,123.5,-125.5</points>
<connection>
<GID>791</GID>
<name>IN_0</name></connection>
<connection>
<GID>793</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1365 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,-136,-42.5,-136</points>
<connection>
<GID>1293</GID>
<name>IN_0</name></connection>
<connection>
<GID>1280</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1015 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127.5,-127.5,127.5,-127.5</points>
<connection>
<GID>792</GID>
<name>IN_0</name></connection>
<connection>
<GID>812</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1271 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-25.5,24,-15.5</points>
<connection>
<GID>1158</GID>
<name>IN_0</name></connection>
<connection>
<GID>1020</GID>
<name>IN_0</name></connection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24,-15.5,41,-15.5</points>
<connection>
<GID>1125</GID>
<name>IN_0</name></connection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>1246 </ID>
<shape>
<vsegment>
<ID>1</ID>
<points>34,-23.5,34,-17.5</points>
<connection>
<GID>1123</GID>
<name>OUT_0</name></connection>
<intersection>-23.5 4</intersection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>34,-17.5,41,-17.5</points>
<connection>
<GID>1125</GID>
<name>IN_1</name></connection>
<intersection>34 1</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>34,-23.5,41,-23.5</points>
<connection>
<GID>1156</GID>
<name>IN_1</name></connection>
<intersection>34 1</intersection></hsegment></shape></wire>
<wire>
<ID>1247 </ID>
<shape>
<vsegment>
<ID>5</ID>
<points>41,-21.5,41,-19.5</points>
<connection>
<GID>1121</GID>
<name>IN_0</name></connection>
<connection>
<GID>1156</GID>
<name>IN_0</name></connection>
<connection>
<GID>1125</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>1014 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127.5,-125.5,127.5,-125.5</points>
<connection>
<GID>793</GID>
<name>OUT_0</name></connection>
<connection>
<GID>812</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1272 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28,-25.5,41,-25.5</points>
<connection>
<GID>1156</GID>
<name>IN_2</name></connection>
<connection>
<GID>1158</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1006 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131.5,-102,132.5,-102</points>
<connection>
<GID>795</GID>
<name>OUT</name></connection>
<connection>
<GID>808</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1357 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46,-109,-46,-109</points>
<connection>
<GID>1269</GID>
<name>IN_1</name></connection>
<connection>
<GID>1270</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1007 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131.5,-104,132.5,-104</points>
<connection>
<GID>808</GID>
<name>IN_1</name></connection>
<intersection>131.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>131.5,-106,131.5,-104</points>
<connection>
<GID>797</GID>
<name>OUT</name></connection>
<intersection>-104 1</intersection></vsegment></shape></wire>
<wire>
<ID>1261 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-128,19,-128</points>
<connection>
<GID>1141</GID>
<name>J</name></connection>
<connection>
<GID>1144</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1262 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-133,19,-132</points>
<connection>
<GID>1146</GID>
<name>OUT</name></connection>
<connection>
<GID>1141</GID>
<name>K</name></connection></vsegment></shape></wire>
<wire>
<ID>1260 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-130,19,-130</points>
<connection>
<GID>1141</GID>
<name>clock</name></connection>
<connection>
<GID>1140</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>95 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161.5,-107.5,161.5,-104</points>
<connection>
<GID>818</GID>
<name>IN_6</name></connection>
<connection>
<GID>818</GID>
<name>IN_4</name></connection>
<connection>
<GID>818</GID>
<name>IN_5</name></connection>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1259 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-128,25,-128</points>
<connection>
<GID>1141</GID>
<name>Q</name></connection>
<connection>
<GID>1142</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1029 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139.5,-123.5,139.5,-123.5</points>
<connection>
<GID>816</GID>
<name>IN_0</name></connection>
<connection>
<GID>826</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>1035 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,-106.5,160,-103</points>
<intersection>-106.5 2</intersection>
<intersection>-103 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>160,-103,161.5,-103</points>
<connection>
<GID>818</GID>
<name>IN_7</name></connection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>145.5,-106.5,160,-106.5</points>
<intersection>145.5 3</intersection>
<intersection>160 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>145.5,-124.5,145.5,-106.5</points>
<connection>
<GID>816</GID>
<name>OUT</name></connection>
<intersection>-106.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>1268 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-133,51,-132</points>
<connection>
<GID>1154</GID>
<name>OUT</name></connection>
<connection>
<GID>1149</GID>
<name>K</name></connection></vsegment></shape></wire>
<wire>
<ID>1290 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-43,-23,-39.5,-23</points>
<connection>
<GID>1178</GID>
<name>IN_0</name></connection>
<connection>
<GID>1181</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1265 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-128,57,-128</points>
<connection>
<GID>1149</GID>
<name>Q</name></connection>
<connection>
<GID>1152</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1031 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160.5,-99,160.5,-95.5</points>
<intersection>-99 1</intersection>
<intersection>-95.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>160.5,-99,161.5,-99</points>
<connection>
<GID>818</GID>
<name>IN_0</name></connection>
<intersection>160.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>146,-95.5,160.5,-95.5</points>
<intersection>146 3</intersection>
<intersection>160.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>146,-95.5,146,-82.5</points>
<intersection>-95.5 2</intersection>
<intersection>-82.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>145.5,-82.5,146,-82.5</points>
<connection>
<GID>820</GID>
<name>OUT</name></connection>
<intersection>146 3</intersection></hsegment></shape></wire>
<wire>
<ID>1058 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159.5,-101,159.5,-96.5</points>
<intersection>-101 1</intersection>
<intersection>-96.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>159.5,-101,161.5,-101</points>
<connection>
<GID>818</GID>
<name>IN_2</name></connection>
<intersection>159.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>145.5,-96.5,159.5,-96.5</points>
<connection>
<GID>864</GID>
<name>OUT</name></connection>
<intersection>159.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1291 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47,-21,-39.5,-21</points>
<connection>
<GID>1176</GID>
<name>IN_1</name></connection>
<intersection>-47 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-47,-23,-47,-21</points>
<connection>
<GID>1181</GID>
<name>IN_0</name></connection>
<connection>
<GID>1165</GID>
<name>IN_0</name></connection>
<intersection>-21 1</intersection></vsegment></shape></wire>
<wire>
<ID>1042 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>180,-87.5,180,-87.5</points>
<connection>
<GID>833</GID>
<name>IN_0</name></connection>
<connection>
<GID>843</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>589 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-54,-62.5,-46.5,-62.5</points>
<connection>
<GID>1234</GID>
<name>IN_0</name></connection>
<connection>
<GID>325</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1263 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-132,13,-132</points>
<connection>
<GID>1147</GID>
<name>IN_0</name></connection>
<connection>
<GID>1146</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1287 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-50.5,-19,-39.5,-19</points>
<connection>
<GID>1176</GID>
<name>IN_0</name></connection>
<intersection>-50.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-50.5,-25,-50.5,-19</points>
<connection>
<GID>1174</GID>
<name>OUT</name></connection>
<intersection>-25 12</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>-50.5,-25,-39.5,-25</points>
<connection>
<GID>1178</GID>
<name>IN_1</name></connection>
<intersection>-50.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>1289 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33.5,-24,-33.5,-24</points>
<connection>
<GID>1178</GID>
<name>OUT</name></connection>
<connection>
<GID>1179</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1050 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113.5,-149,113.5,-149</points>
<connection>
<GID>848</GID>
<name>IN_0</name></connection>
<connection>
<GID>857</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>1047 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100.5,-145,100.5,-145</points>
<connection>
<GID>850</GID>
<name>IN_0</name></connection>
<connection>
<GID>855</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1167 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-36,18,-36</points>
<connection>
<GID>1027</GID>
<name>IN_0</name></connection>
<connection>
<GID>1039</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1048 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100.5,-147,100.5,-147</points>
<connection>
<GID>851</GID>
<name>IN_0</name></connection>
<connection>
<GID>855</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1157 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244.5,-67,244.5,-52.5</points>
<intersection>-67 2</intersection>
<intersection>-52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>244.5,-52.5,258.5,-52.5</points>
<connection>
<GID>1011</GID>
<name>IN_7</name></connection>
<intersection>244.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>243.5,-67,244.5,-67</points>
<connection>
<GID>994</GID>
<name>IN_0</name></connection>
<intersection>244.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>353 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-61,27.5,-60</points>
<intersection>-61 1</intersection>
<intersection>-60 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-61,31.5,-61</points>
<connection>
<GID>249</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-60,27.5,-60</points>
<connection>
<GID>1084</GID>
<name>OUT</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1046 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>100.5,-149,100.5,-149</points>
<connection>
<GID>852</GID>
<name>IN_0</name></connection>
<connection>
<GID>855</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1049 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100.5,-151,100.5,-151</points>
<connection>
<GID>853</GID>
<name>IN_0</name></connection>
<connection>
<GID>855</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>1170 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-46,18,-46</points>
<connection>
<GID>1040</GID>
<name>IN_2</name></connection>
<intersection>-46 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-46,18,-46</points>
<connection>
<GID>1032</GID>
<name>IN_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>1052 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>107.5,-148,107.5,-148</points>
<connection>
<GID>855</GID>
<name>OUT</name></connection>
<connection>
<GID>857</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1051 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-153,107.5,-150</points>
<connection>
<GID>857</GID>
<name>IN_1</name></connection>
<intersection>-153 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100.5,-153,107.5,-153</points>
<connection>
<GID>858</GID>
<name>IN_0</name></connection>
<intersection>107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1174 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-48,18,-48</points>
<connection>
<GID>1035</GID>
<name>IN_0</name></connection>
<connection>
<GID>1041</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1055 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134.5,-149,134.5,-149</points>
<connection>
<GID>859</GID>
<name>IN_0</name></connection>
<connection>
<GID>862</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>1053 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128.5,-148,128.5,-148</points>
<connection>
<GID>860</GID>
<name>IN_0</name></connection>
<connection>
<GID>862</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>361 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-54,-37,-46.5,-37</points>
<connection>
<GID>1197</GID>
<name>IN_0</name></connection>
<connection>
<GID>275</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1054 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128.5,-150,128.5,-150</points>
<connection>
<GID>861</GID>
<name>IN_0</name></connection>
<connection>
<GID>862</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1171 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-42,18,-42</points>
<connection>
<GID>1040</GID>
<name>IN_0</name></connection>
<connection>
<GID>1031</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1177 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24,-44,33,-44</points>
<connection>
<GID>1040</GID>
<name>OUT</name></connection>
<connection>
<GID>1043</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1059 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>139.5,-94.5,139.5,-94.5</points>
<connection>
<GID>864</GID>
<name>IN_0</name></connection>
<connection>
<GID>865</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1060 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169,-149,169,-149</points>
<connection>
<GID>866</GID>
<name>IN_0</name></connection>
<connection>
<GID>872</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>1176 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>24,-42,33,-42</points>
<connection>
<GID>1043</GID>
<name>IN_0</name></connection>
<intersection>24 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>24,-42,24,-38</points>
<connection>
<GID>1039</GID>
<name>OUT</name></connection>
<intersection>-42 2</intersection></vsegment></shape></wire>
<wire>
<ID>1178 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>24,-46,33,-46</points>
<connection>
<GID>1043</GID>
<name>IN_2</name></connection>
<intersection>24 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>24,-50,24,-46</points>
<connection>
<GID>1041</GID>
<name>OUT</name></connection>
<intersection>-46 2</intersection></vsegment></shape></wire>
<wire>
<ID>1064 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157,-151,157,-151</points>
<connection>
<GID>867</GID>
<name>IN_0</name></connection>
<connection>
<GID>875</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1065 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157,-153,157,-153</points>
<connection>
<GID>868</GID>
<name>IN_0</name></connection>
<connection>
<GID>875</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>576 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>252.5,-28.5,252.5,-26.5</points>
<connection>
<GID>346</GID>
<name>IN_1</name></connection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>252.5,-28.5,252.5,-28.5</points>
<connection>
<GID>284</GID>
<name>OUT_0</name></connection>
<intersection>252.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1062 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>155,-145,157,-145</points>
<connection>
<GID>869</GID>
<name>IN_0</name></connection>
<connection>
<GID>874</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1063 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>155,-147,157,-147</points>
<connection>
<GID>870</GID>
<name>IN_0</name></connection>
<connection>
<GID>874</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1073 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-173,121.5,-173</points>
<connection>
<GID>877</GID>
<name>IN_0</name></connection>
<connection>
<GID>881</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>1191 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-48.5,43,-48.5</points>
<connection>
<GID>1056</GID>
<name>IN_0</name></connection>
<connection>
<GID>1052</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1194 </ID>
<shape>
<hsegment>
<ID>9</ID>
<points>49,-48,50,-48</points>
<connection>
<GID>1037</GID>
<name>K</name></connection>
<intersection>49 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>49,-49.5,49,-48</points>
<connection>
<GID>1056</GID>
<name>OUT</name></connection>
<intersection>-48 9</intersection></vsegment></shape></wire>
<wire>
<ID>1072 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-172,115.5,-172</points>
<connection>
<GID>879</GID>
<name>OUT_0</name></connection>
<connection>
<GID>881</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1071 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-174,115.5,-174</points>
<connection>
<GID>880</GID>
<name>IN_0</name></connection>
<connection>
<GID>881</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1075 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145.5,-174,145.5,-174</points>
<connection>
<GID>884</GID>
<name>IN_0</name></connection>
<connection>
<GID>885</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1077 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151.5,-173,151.5,-173</points>
<connection>
<GID>885</GID>
<name>OUT</name></connection>
<connection>
<GID>886</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1198 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-81.5,22.5,-81.5</points>
<connection>
<GID>1064</GID>
<name>IN_0</name></connection>
<connection>
<GID>1068</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1211 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-63,18,-63</points>
<connection>
<GID>1093</GID>
<name>IN_0</name></connection>
<connection>
<GID>1086</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1081 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-193,121.5,-193</points>
<connection>
<GID>889</GID>
<name>IN_0</name></connection>
<connection>
<GID>893</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>1079 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-194,115.5,-194</points>
<connection>
<GID>892</GID>
<name>IN_0</name></connection>
<connection>
<GID>893</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1222 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-87.5,27.5,-84.5</points>
<intersection>-87.5 2</intersection>
<intersection>-84.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-84.5,29,-84.5</points>
<connection>
<GID>1096</GID>
<name>IN_3</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-87.5,27.5,-87.5</points>
<connection>
<GID>1072</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1087 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145.5,-192,145.5,-192</points>
<connection>
<GID>894</GID>
<name>IN_0</name></connection>
<connection>
<GID>896</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1085 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151.5,-193,151.5,-193</points>
<connection>
<GID>896</GID>
<name>OUT</name></connection>
<connection>
<GID>897</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1088 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-202,84,-202</points>
<connection>
<GID>901</GID>
<name>IN_0</name></connection>
<connection>
<GID>916</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1089 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-204,84,-204</points>
<connection>
<GID>902</GID>
<name>IN_0</name></connection>
<connection>
<GID>916</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1092 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-208.5,90,-206.5</points>
<connection>
<GID>918</GID>
<name>IN_1</name></connection>
<intersection>-208.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>84,-208.5,90,-208.5</points>
<connection>
<GID>904</GID>
<name>IN_0</name></connection>
<intersection>90 0</intersection></hsegment></shape></wire>
<wire>
<ID>1090 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-206,84,-206</points>
<connection>
<GID>905</GID>
<name>IN_0</name></connection>
<connection>
<GID>916</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>382 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46.5,-48,-46.5,-48</points>
<connection>
<GID>1208</GID>
<name>IN_0</name></connection>
<connection>
<GID>287</GID>
<name>IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>1097 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-218,90,-215.5</points>
<connection>
<GID>922</GID>
<name>IN_1</name></connection>
<intersection>-218 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>84,-218,90,-218</points>
<connection>
<GID>907</GID>
<name>IN_0</name></connection>
<intersection>90 0</intersection></hsegment></shape></wire>
<wire>
<ID>1345 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40,-86,-40,-86</points>
<connection>
<GID>1242</GID>
<name>IN_0</name></connection>
<connection>
<GID>1253</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>1095 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-215.5,84,-215.5</points>
<connection>
<GID>908</GID>
<name>IN_0</name></connection>
<connection>
<GID>920</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>1018 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-39.5,-63,-39.5,-60</points>
<connection>
<GID>1190</GID>
<name>IN_1</name></connection>
<connection>
<GID>325</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>1195 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-46,50,-46</points>
<connection>
<GID>1057</GID>
<name>IN_0</name></connection>
<connection>
<GID>1037</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>1094 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-213.5,84,-213.5</points>
<connection>
<GID>910</GID>
<name>IN_0</name></connection>
<connection>
<GID>920</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1093 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-211.5,84,-211.5</points>
<connection>
<GID>912</GID>
<name>IN_0</name></connection>
<connection>
<GID>920</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1099 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-221.5,90,-221.5</points>
<connection>
<GID>913</GID>
<name>IN_0</name></connection>
<connection>
<GID>924</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1098 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-223.5,90,-223.5</points>
<connection>
<GID>914</GID>
<name>IN_0</name></connection>
<connection>
<GID>924</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1209 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-61,18,-61</points>
<connection>
<GID>1091</GID>
<name>IN_0</name></connection>
<connection>
<GID>1084</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1091 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-204.5,90,-204</points>
<connection>
<GID>918</GID>
<name>IN_0</name></connection>
<connection>
<GID>916</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>1196 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-85,52.5,-85</points>
<connection>
<GID>1058</GID>
<name>Q</name></connection>
<connection>
<GID>1060</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>16 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96,-212.5,96,-205.5</points>
<connection>
<GID>918</GID>
<name>OUT</name></connection>
<connection>
<GID>926</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1096 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-213.5,90,-213.5</points>
<connection>
<GID>920</GID>
<name>OUT</name></connection>
<connection>
<GID>922</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1343 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46,-85,-46,-85</points>
<connection>
<GID>1253</GID>
<name>IN_0</name></connection>
<connection>
<GID>1254</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1100 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>96,-214.5,96,-214.5</points>
<connection>
<GID>922</GID>
<name>OUT</name></connection>
<connection>
<GID>926</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1105 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,-213,120,-213</points>
<connection>
<GID>929</GID>
<name>IN_0</name></connection>
<connection>
<GID>930</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1106 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,-215,120,-215</points>
<connection>
<GID>929</GID>
<name>IN_1</name></connection>
<connection>
<GID>931</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1356 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46,-107,-46,-107</points>
<connection>
<GID>1269</GID>
<name>IN_0</name></connection>
<connection>
<GID>1267</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1355 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40,-108,-40,-108</points>
<connection>
<GID>1269</GID>
<name>OUT</name></connection>
<connection>
<GID>1246</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>752 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-54,-66.5,-46.5,-66.5</points>
<connection>
<GID>325</GID>
<name>IN_4</name></connection>
<connection>
<GID>1238</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1110 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187.5,-215,187.5,-215</points>
<connection>
<GID>938</GID>
<name>IN_0</name></connection>
<connection>
<GID>940</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>431 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-54,-58.5,-46.5,-58.5</points>
<connection>
<GID>1230</GID>
<name>IN_0</name></connection>
<connection>
<GID>313</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1116 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181.5,-214,181.5,-213</points>
<connection>
<GID>948</GID>
<name>OUT</name></connection>
<connection>
<GID>940</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1113 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181.5,-217,181.5,-216</points>
<connection>
<GID>943</GID>
<name>OUT</name></connection>
<connection>
<GID>940</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1245 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-20.5,30,-20.5</points>
<connection>
<GID>1120</GID>
<name>IN_0</name></connection>
<connection>
<GID>1123</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1115 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>175.5,-212,175.5,-212</points>
<connection>
<GID>946</GID>
<name>IN_0</name></connection>
<connection>
<GID>948</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1270 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-134,45,-134</points>
<connection>
<GID>1154</GID>
<name>IN_1</name></connection>
<connection>
<GID>1155</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1119 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-108.5,-41,-108.5,-41</points>
<connection>
<GID>951</GID>
<name>IN_0</name></connection>
<connection>
<GID>954</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>1118 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-114.5,-40,-114.5,-40</points>
<connection>
<GID>952</GID>
<name>IN_0</name></connection>
<connection>
<GID>954</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1117 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-114.5,-42,-114.5,-42</points>
<connection>
<GID>953</GID>
<name>IN_0</name></connection>
<connection>
<GID>954</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1129 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228.5,-24.5,228.5,-24.5</points>
<connection>
<GID>959</GID>
<name>IN_0</name></connection>
<connection>
<GID>969</GID>
<name>OUT_2</name></connection></vsegment></shape></wire>
<wire>
<ID>1127 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228.5,-26.5,228.5,-26.5</points>
<connection>
<GID>961</GID>
<name>IN_0</name></connection>
<connection>
<GID>969</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1363 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,-132,-42.5,-132</points>
<connection>
<GID>1291</GID>
<name>IN_0</name></connection>
<connection>
<GID>1278</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1128 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>228.5,-25.5,233.5,-25.5</points>
<connection>
<GID>962</GID>
<name>IN_0</name></connection>
<connection>
<GID>969</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1372 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,-150,-42.5,-150</points>
<connection>
<GID>1300</GID>
<name>IN_0</name></connection>
<connection>
<GID>1287</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1130 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>228.5,-23.5,233.5,-23.5</points>
<connection>
<GID>963</GID>
<name>IN_0</name></connection>
<connection>
<GID>969</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1132 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>228.5,-21.5,233.5,-21.5</points>
<connection>
<GID>965</GID>
<name>IN_0</name></connection>
<connection>
<GID>969</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1212 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-65,18,-65</points>
<connection>
<GID>1086</GID>
<name>IN_1</name></connection>
<connection>
<GID>1094</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1152 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>265.5,-52,265.5,-52</points>
<connection>
<GID>973</GID>
<name>IN_0</name></connection>
<connection>
<GID>1011</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>1148 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>237.5,-43,237.5,-43</points>
<connection>
<GID>977</GID>
<name>IN_0</name></connection>
<connection>
<GID>1007</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1139 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230.5,-47.5,230.5,-47.5</points>
<connection>
<GID>982</GID>
<name>IN_0</name></connection>
<connection>
<GID>997</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1137 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230.5,-49.5,230.5,-49.5</points>
<connection>
<GID>984</GID>
<name>IN_0</name></connection>
<connection>
<GID>997</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>1143 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>237.5,-53.5,237.5,-50.5</points>
<connection>
<GID>999</GID>
<name>IN_1</name></connection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>230.5,-53.5,237.5,-53.5</points>
<connection>
<GID>990</GID>
<name>IN_0</name></connection>
<intersection>237.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1150 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>237.5,-62.5,237.5,-62.5</points>
<connection>
<GID>992</GID>
<name>IN_0</name></connection>
<connection>
<GID>1009</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1151 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>237.5,-64.5,237.5,-64.5</points>
<connection>
<GID>993</GID>
<name>IN_0</name></connection>
<connection>
<GID>1009</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1284 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33.5,-20,-33.5,-20</points>
<connection>
<GID>1176</GID>
<name>OUT</name></connection>
<connection>
<GID>1161</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1154 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>243.5,-49.5,258.5,-49.5</points>
<connection>
<GID>999</GID>
<name>OUT</name></connection>
<connection>
<GID>1011</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1156 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244,-63.5,244,-51.5</points>
<intersection>-63.5 2</intersection>
<intersection>-51.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>244,-51.5,258.5,-51.5</points>
<connection>
<GID>1011</GID>
<name>IN_3</name></connection>
<intersection>244 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>243.5,-63.5,244,-63.5</points>
<connection>
<GID>1009</GID>
<name>OUT</name></connection>
<intersection>244 0</intersection></hsegment></shape></wire>
<wire>
<ID>587 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>245.5,-54.5,258.5,-54.5</points>
<connection>
<GID>1011</GID>
<name>IN_5</name></connection>
<intersection>245.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>245.5,-71,245.5,-54.5</points>
<intersection>-71 4</intersection>
<intersection>-54.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>243.5,-71,245.5,-71</points>
<connection>
<GID>375</GID>
<name>IN_0</name></connection>
<intersection>245.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>1165 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-44,56,-44</points>
<connection>
<GID>1025</GID>
<name>IN_0</name></connection>
<connection>
<GID>1037</GID>
<name>Q</name></connection></vsegment></shape></wire>
<wire>
<ID>1168 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-40,18,-40</points>
<connection>
<GID>1029</GID>
<name>IN_0</name></connection>
<connection>
<GID>1039</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>344 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126,-218.5,126,-216</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<connection>
<GID>147</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1213 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35,-85,46.5,-85</points>
<connection>
<GID>1096</GID>
<name>OUT</name></connection>
<connection>
<GID>1058</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>1219 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-81.5,29,-81.5</points>
<connection>
<GID>1096</GID>
<name>IN_0</name></connection>
<connection>
<GID>1068</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>358 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46.5,-36,-46.5,-36</points>
<connection>
<GID>275</GID>
<name>IN_2</name></connection>
<connection>
<GID>1196</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1201 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-90,20.5,-90</points>
<connection>
<GID>1076</GID>
<name>IN_0</name></connection>
<connection>
<GID>1078</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1208 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-55,18,-55</points>
<connection>
<GID>1082</GID>
<name>IN_0</name></connection>
<connection>
<GID>1088</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>356 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46.5,-38,-46.5,-38</points>
<connection>
<GID>275</GID>
<name>IN_7</name></connection>
<connection>
<GID>1198</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1207 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-57,18,-57</points>
<connection>
<GID>1082</GID>
<name>IN_1</name></connection>
<connection>
<GID>1087</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1210 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-59,18,-59</points>
<connection>
<GID>1084</GID>
<name>IN_0</name></connection>
<connection>
<GID>1092</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1229 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-110,43,-110</points>
<connection>
<GID>1102</GID>
<name>IN_0</name></connection>
<connection>
<GID>1103</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>1228 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-108,49,-108</points>
<connection>
<GID>1103</GID>
<name>Q</name></connection>
<connection>
<GID>1104</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>598 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-54,-64.5,-46.5,-64.5</points>
<connection>
<GID>325</GID>
<name>IN_6</name></connection>
<connection>
<GID>1236</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1264 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-134,13,-134</points>
<connection>
<GID>1146</GID>
<name>IN_1</name></connection>
<connection>
<GID>1148</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>569 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>263,-39,263,-39</points>
<connection>
<GID>335</GID>
<name>IN_0</name></connection>
<connection>
<GID>322</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1283 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-56.5,-21,-56.5,-21</points>
<connection>
<GID>1164</GID>
<name>IN_0</name></connection>
<connection>
<GID>1174</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1299 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33.5,-59,-33.5,-59</points>
<connection>
<GID>1190</GID>
<name>OUT</name></connection>
<connection>
<GID>1193</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1346 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-46,-90.5,-40,-90.5</points>
<connection>
<GID>1243</GID>
<name>IN_0</name></connection>
<connection>
<GID>1256</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1364 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,-134,-42.5,-134</points>
<connection>
<GID>1292</GID>
<name>IN_0</name></connection>
<connection>
<GID>1279</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1350 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52,-99.5,-52,-99.5</points>
<connection>
<GID>1261</GID>
<name>IN_0</name></connection>
<connection>
<GID>1262</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1353 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46,-100.5,-46,-100.5</points>
<connection>
<GID>1261</GID>
<name>OUT</name></connection>
<connection>
<GID>1265</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1362 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,-130,-42.5,-130</points>
<connection>
<GID>1290</GID>
<name>IN_0</name></connection>
<connection>
<GID>1277</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>349 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-67,18,-67</points>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<connection>
<GID>39</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>350 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-69,18,-69</points>
<connection>
<GID>245</GID>
<name>IN_0</name></connection>
<connection>
<GID>39</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>351 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-62,38.5,-50.5</points>
<connection>
<GID>249</GID>
<name>OUT</name></connection>
<intersection>-50.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>38.5,-50.5,43,-50.5</points>
<connection>
<GID>1056</GID>
<name>IN_1</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>352 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-59,27.5,-56</points>
<intersection>-59 1</intersection>
<intersection>-56 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-59,31.5,-59</points>
<connection>
<GID>249</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-56,27.5,-56</points>
<connection>
<GID>1082</GID>
<name>OUT</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>354 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-64,27.5,-63</points>
<intersection>-64 2</intersection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-63,31.5,-63</points>
<connection>
<GID>249</GID>
<name>IN_2</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-64,27.5,-64</points>
<connection>
<GID>1086</GID>
<name>OUT</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>360 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-54,-35,-46.5,-35</points>
<connection>
<GID>275</GID>
<name>IN_1</name></connection>
<connection>
<GID>1195</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>362 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-54,-39,-46.5,-39</points>
<connection>
<GID>275</GID>
<name>IN_6</name></connection>
<connection>
<GID>1199</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>363 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-54,-41,-46.5,-41</points>
<connection>
<GID>1201</GID>
<name>IN_0</name></connection>
<connection>
<GID>275</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>381 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46.5,-44,-46.5,-44</points>
<connection>
<GID>1204</GID>
<name>IN_0</name></connection>
<connection>
<GID>287</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>384 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46.5,-46,-46.5,-46</points>
<connection>
<GID>1206</GID>
<name>IN_0</name></connection>
<connection>
<GID>287</GID>
<name>IN_7</name></connection></vsegment></shape></wire>
<wire>
<ID>386 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-54,-45,-46.5,-45</points>
<connection>
<GID>287</GID>
<name>IN_3</name></connection>
<connection>
<GID>1205</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>387 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-54,-47,-46.5,-47</points>
<connection>
<GID>1207</GID>
<name>IN_0</name></connection>
<connection>
<GID>287</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>389 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-39.5,-45.5,-39.5,-42.5</points>
<connection>
<GID>1188</GID>
<name>IN_1</name></connection>
<connection>
<GID>287</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>391 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46.5,-51.5,-46.5,-51.5</points>
<connection>
<GID>1210</GID>
<name>IN_0</name></connection>
<connection>
<GID>313</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>392 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46.5,-53.5,-46.5,-53.5</points>
<connection>
<GID>1225</GID>
<name>IN_0</name></connection>
<connection>
<GID>313</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>394 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-54,-52.5,-46.5,-52.5</points>
<connection>
<GID>313</GID>
<name>IN_1</name></connection>
<connection>
<GID>1224</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>395 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-54,-54.5,-46.5,-54.5</points>
<connection>
<GID>1226</GID>
<name>IN_0</name></connection>
<connection>
<GID>313</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>538 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46.5,-59.5,-46.5,-59.5</points>
<connection>
<GID>325</GID>
<name>IN_0</name></connection>
<connection>
<GID>1231</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>552 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46.5,-63.5,-46.5,-63.5</points>
<connection>
<GID>325</GID>
<name>IN_7</name></connection>
<connection>
<GID>1235</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>562 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46.5,-65.5,-46.5,-65.5</points>
<connection>
<GID>325</GID>
<name>IN_5</name></connection>
<connection>
<GID>1237</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>567 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-54,-60.5,-46.5,-60.5</points>
<connection>
<GID>325</GID>
<name>IN_1</name></connection>
<connection>
<GID>1232</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1017 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-39.5,-58,-39.5,-55</points>
<connection>
<GID>1190</GID>
<name>IN_0</name></connection>
<connection>
<GID>313</GID>
<name>OUT</name></connection></vsegment></shape></wire></page 2></circuit>